// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     Jun 12 2021 20:10:07

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    led,
    usb_tx,
    usb_rx,
    rst_n,
    clk);

    output [7:0] led;
    output usb_tx;
    input usb_rx;
    input rst_n;
    input clk;

    wire N__3165;
    wire N__3164;
    wire N__3163;
    wire N__3154;
    wire N__3153;
    wire N__3152;
    wire N__3145;
    wire N__3144;
    wire N__3143;
    wire N__3136;
    wire N__3135;
    wire N__3134;
    wire N__3127;
    wire N__3126;
    wire N__3125;
    wire N__3118;
    wire N__3117;
    wire N__3116;
    wire N__3109;
    wire N__3108;
    wire N__3107;
    wire N__3100;
    wire N__3099;
    wire N__3098;
    wire N__3091;
    wire N__3090;
    wire N__3089;
    wire N__3082;
    wire N__3081;
    wire N__3080;
    wire N__3073;
    wire N__3072;
    wire N__3071;
    wire N__3064;
    wire N__3063;
    wire N__3062;
    wire N__3045;
    wire N__3044;
    wire N__3041;
    wire N__3038;
    wire N__3033;
    wire N__3032;
    wire N__3029;
    wire N__3026;
    wire N__3021;
    wire N__3018;
    wire N__3017;
    wire N__3014;
    wire N__3011;
    wire N__3006;
    wire N__3003;
    wire N__3000;
    wire N__2997;
    wire N__2996;
    wire N__2993;
    wire N__2990;
    wire N__2985;
    wire N__2984;
    wire N__2981;
    wire N__2978;
    wire N__2977;
    wire N__2976;
    wire N__2975;
    wire N__2974;
    wire N__2973;
    wire N__2972;
    wire N__2969;
    wire N__2966;
    wire N__2965;
    wire N__2964;
    wire N__2961;
    wire N__2960;
    wire N__2959;
    wire N__2954;
    wire N__2947;
    wire N__2944;
    wire N__2941;
    wire N__2940;
    wire N__2939;
    wire N__2934;
    wire N__2931;
    wire N__2926;
    wire N__2921;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2895;
    wire N__2892;
    wire N__2889;
    wire N__2888;
    wire N__2887;
    wire N__2886;
    wire N__2885;
    wire N__2884;
    wire N__2881;
    wire N__2880;
    wire N__2879;
    wire N__2878;
    wire N__2877;
    wire N__2876;
    wire N__2875;
    wire N__2874;
    wire N__2873;
    wire N__2872;
    wire N__2871;
    wire N__2870;
    wire N__2865;
    wire N__2860;
    wire N__2859;
    wire N__2858;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2842;
    wire N__2837;
    wire N__2832;
    wire N__2825;
    wire N__2820;
    wire N__2817;
    wire N__2812;
    wire N__2809;
    wire N__2790;
    wire N__2789;
    wire N__2786;
    wire N__2783;
    wire N__2778;
    wire N__2777;
    wire N__2776;
    wire N__2775;
    wire N__2774;
    wire N__2773;
    wire N__2772;
    wire N__2771;
    wire N__2768;
    wire N__2765;
    wire N__2764;
    wire N__2757;
    wire N__2750;
    wire N__2743;
    wire N__2740;
    wire N__2733;
    wire N__2732;
    wire N__2729;
    wire N__2728;
    wire N__2727;
    wire N__2726;
    wire N__2725;
    wire N__2724;
    wire N__2723;
    wire N__2722;
    wire N__2715;
    wire N__2708;
    wire N__2701;
    wire N__2694;
    wire N__2693;
    wire N__2692;
    wire N__2691;
    wire N__2690;
    wire N__2689;
    wire N__2686;
    wire N__2685;
    wire N__2684;
    wire N__2683;
    wire N__2680;
    wire N__2677;
    wire N__2674;
    wire N__2671;
    wire N__2664;
    wire N__2657;
    wire N__2650;
    wire N__2643;
    wire N__2642;
    wire N__2641;
    wire N__2640;
    wire N__2639;
    wire N__2638;
    wire N__2637;
    wire N__2636;
    wire N__2635;
    wire N__2632;
    wire N__2627;
    wire N__2620;
    wire N__2613;
    wire N__2604;
    wire N__2601;
    wire N__2598;
    wire N__2595;
    wire N__2592;
    wire N__2589;
    wire N__2588;
    wire N__2585;
    wire N__2584;
    wire N__2581;
    wire N__2578;
    wire N__2575;
    wire N__2572;
    wire N__2569;
    wire N__2566;
    wire N__2563;
    wire N__2558;
    wire N__2553;
    wire N__2552;
    wire N__2551;
    wire N__2550;
    wire N__2549;
    wire N__2548;
    wire N__2547;
    wire N__2546;
    wire N__2545;
    wire N__2544;
    wire N__2543;
    wire N__2542;
    wire N__2541;
    wire N__2540;
    wire N__2539;
    wire N__2508;
    wire N__2505;
    wire N__2502;
    wire N__2499;
    wire N__2498;
    wire N__2495;
    wire N__2492;
    wire N__2489;
    wire N__2484;
    wire N__2483;
    wire N__2480;
    wire N__2477;
    wire N__2474;
    wire N__2469;
    wire N__2468;
    wire N__2465;
    wire N__2462;
    wire N__2457;
    wire N__2454;
    wire N__2451;
    wire N__2450;
    wire N__2447;
    wire N__2444;
    wire N__2439;
    wire N__2438;
    wire N__2435;
    wire N__2432;
    wire N__2427;
    wire N__2426;
    wire N__2423;
    wire N__2420;
    wire N__2415;
    wire N__2412;
    wire N__2411;
    wire N__2408;
    wire N__2405;
    wire N__2400;
    wire N__2397;
    wire N__2396;
    wire N__2393;
    wire N__2390;
    wire N__2385;
    wire N__2382;
    wire N__2379;
    wire N__2376;
    wire N__2373;
    wire N__2370;
    wire N__2367;
    wire N__2364;
    wire N__2363;
    wire N__2362;
    wire N__2355;
    wire N__2352;
    wire N__2351;
    wire N__2348;
    wire N__2347;
    wire N__2346;
    wire N__2339;
    wire N__2336;
    wire N__2331;
    wire N__2330;
    wire N__2329;
    wire N__2328;
    wire N__2325;
    wire N__2322;
    wire N__2319;
    wire N__2316;
    wire N__2307;
    wire N__2306;
    wire N__2303;
    wire N__2300;
    wire N__2295;
    wire N__2292;
    wire N__2289;
    wire N__2286;
    wire N__2283;
    wire N__2280;
    wire N__2277;
    wire N__2274;
    wire N__2271;
    wire N__2268;
    wire N__2267;
    wire N__2266;
    wire N__2265;
    wire N__2264;
    wire N__2261;
    wire N__2258;
    wire N__2255;
    wire N__2250;
    wire N__2241;
    wire N__2238;
    wire N__2235;
    wire N__2232;
    wire N__2229;
    wire N__2228;
    wire N__2227;
    wire N__2226;
    wire N__2223;
    wire N__2220;
    wire N__2217;
    wire N__2216;
    wire N__2213;
    wire N__2212;
    wire N__2209;
    wire N__2208;
    wire N__2207;
    wire N__2204;
    wire N__2201;
    wire N__2198;
    wire N__2193;
    wire N__2190;
    wire N__2185;
    wire N__2172;
    wire N__2171;
    wire N__2170;
    wire N__2169;
    wire N__2166;
    wire N__2163;
    wire N__2160;
    wire N__2157;
    wire N__2148;
    wire N__2147;
    wire N__2144;
    wire N__2141;
    wire N__2140;
    wire N__2139;
    wire N__2138;
    wire N__2135;
    wire N__2132;
    wire N__2129;
    wire N__2124;
    wire N__2117;
    wire N__2114;
    wire N__2109;
    wire N__2106;
    wire N__2103;
    wire N__2100;
    wire N__2099;
    wire N__2096;
    wire N__2095;
    wire N__2094;
    wire N__2093;
    wire N__2092;
    wire N__2091;
    wire N__2090;
    wire N__2087;
    wire N__2084;
    wire N__2081;
    wire N__2076;
    wire N__2073;
    wire N__2070;
    wire N__2067;
    wire N__2062;
    wire N__2057;
    wire N__2046;
    wire N__2043;
    wire N__2040;
    wire N__2039;
    wire N__2038;
    wire N__2037;
    wire N__2036;
    wire N__2035;
    wire N__2034;
    wire N__2029;
    wire N__2026;
    wire N__2021;
    wire N__2016;
    wire N__2007;
    wire N__2004;
    wire N__2003;
    wire N__2002;
    wire N__1999;
    wire N__1998;
    wire N__1995;
    wire N__1992;
    wire N__1989;
    wire N__1986;
    wire N__1981;
    wire N__1976;
    wire N__1971;
    wire N__1968;
    wire N__1965;
    wire N__1964;
    wire N__1961;
    wire N__1958;
    wire N__1955;
    wire N__1950;
    wire N__1947;
    wire N__1944;
    wire N__1943;
    wire N__1942;
    wire N__1937;
    wire N__1934;
    wire N__1929;
    wire N__1926;
    wire N__1923;
    wire N__1922;
    wire N__1917;
    wire N__1914;
    wire N__1911;
    wire N__1908;
    wire N__1905;
    wire N__1904;
    wire N__1903;
    wire N__1900;
    wire N__1897;
    wire N__1896;
    wire N__1895;
    wire N__1894;
    wire N__1891;
    wire N__1890;
    wire N__1887;
    wire N__1882;
    wire N__1873;
    wire N__1866;
    wire N__1863;
    wire N__1860;
    wire N__1857;
    wire N__1854;
    wire N__1853;
    wire N__1852;
    wire N__1851;
    wire N__1848;
    wire N__1845;
    wire N__1840;
    wire N__1833;
    wire N__1832;
    wire N__1829;
    wire N__1826;
    wire N__1825;
    wire N__1824;
    wire N__1823;
    wire N__1822;
    wire N__1821;
    wire N__1820;
    wire N__1819;
    wire N__1816;
    wire N__1813;
    wire N__1810;
    wire N__1805;
    wire N__1802;
    wire N__1795;
    wire N__1782;
    wire N__1781;
    wire N__1776;
    wire N__1773;
    wire N__1770;
    wire N__1767;
    wire N__1766;
    wire N__1765;
    wire N__1764;
    wire N__1763;
    wire N__1762;
    wire N__1759;
    wire N__1756;
    wire N__1753;
    wire N__1746;
    wire N__1737;
    wire N__1734;
    wire N__1731;
    wire N__1728;
    wire N__1725;
    wire N__1722;
    wire N__1721;
    wire N__1718;
    wire N__1715;
    wire N__1710;
    wire N__1707;
    wire N__1706;
    wire N__1705;
    wire N__1702;
    wire N__1699;
    wire N__1696;
    wire N__1689;
    wire N__1688;
    wire N__1687;
    wire N__1682;
    wire N__1679;
    wire N__1674;
    wire N__1671;
    wire N__1670;
    wire N__1669;
    wire N__1668;
    wire N__1665;
    wire N__1660;
    wire N__1657;
    wire N__1654;
    wire N__1647;
    wire N__1646;
    wire N__1645;
    wire N__1642;
    wire N__1637;
    wire N__1632;
    wire N__1629;
    wire N__1626;
    wire N__1623;
    wire N__1622;
    wire N__1619;
    wire N__1616;
    wire N__1615;
    wire N__1612;
    wire N__1607;
    wire N__1602;
    wire N__1599;
    wire N__1598;
    wire N__1597;
    wire N__1596;
    wire N__1593;
    wire N__1590;
    wire N__1587;
    wire N__1584;
    wire N__1575;
    wire N__1572;
    wire N__1571;
    wire N__1570;
    wire N__1569;
    wire N__1568;
    wire N__1563;
    wire N__1556;
    wire N__1551;
    wire N__1548;
    wire N__1545;
    wire N__1542;
    wire N__1539;
    wire N__1536;
    wire N__1533;
    wire N__1530;
    wire N__1529;
    wire N__1526;
    wire N__1523;
    wire N__1518;
    wire N__1517;
    wire N__1514;
    wire N__1511;
    wire N__1506;
    wire N__1503;
    wire N__1502;
    wire N__1499;
    wire N__1496;
    wire N__1491;
    wire N__1488;
    wire N__1485;
    wire N__1482;
    wire N__1479;
    wire N__1478;
    wire N__1475;
    wire N__1472;
    wire N__1469;
    wire N__1464;
    wire N__1461;
    wire N__1458;
    wire N__1455;
    wire N__1452;
    wire N__1449;
    wire N__1448;
    wire N__1447;
    wire N__1446;
    wire N__1439;
    wire N__1436;
    wire N__1431;
    wire N__1428;
    wire N__1425;
    wire N__1422;
    wire N__1421;
    wire N__1418;
    wire N__1415;
    wire N__1412;
    wire N__1407;
    wire N__1406;
    wire N__1403;
    wire N__1400;
    wire N__1395;
    wire N__1394;
    wire N__1391;
    wire N__1388;
    wire N__1383;
    wire N__1380;
    wire N__1377;
    wire N__1374;
    wire N__1373;
    wire N__1370;
    wire N__1365;
    wire N__1362;
    wire N__1361;
    wire N__1360;
    wire N__1359;
    wire N__1358;
    wire N__1357;
    wire N__1344;
    wire N__1341;
    wire N__1338;
    wire N__1335;
    wire N__1332;
    wire N__1329;
    wire N__1326;
    wire N__1323;
    wire N__1322;
    wire N__1321;
    wire N__1320;
    wire N__1311;
    wire N__1308;
    wire N__1305;
    wire N__1302;
    wire N__1299;
    wire N__1296;
    wire VCCG0;
    wire GNDG0;
    wire \reset_cond.M_stage_qZ0Z_1 ;
    wire \reset_cond.M_stage_qZ0Z_2 ;
    wire rst_n_c;
    wire \reset_cond.M_stage_qZ0Z_0 ;
    wire \uart_rx.un1_M_ctr_q_5_ac0_5_s_0_0_cascade_ ;
    wire \uart_rx.N_102_0_cascade_ ;
    wire \uart_rx.un1_M_ctr_q_5_ac0_7_0 ;
    wire \uart_rx.N_102_0 ;
    wire \uart_rx.un1_M_ctr_q_5_ac0_5_s_0_0 ;
    wire \uart_tx.M_state_q_ns_0_o2_4_0_cascade_ ;
    wire \uart_tx.N_183_0_cascade_ ;
    wire \uart_tx.M_state_q_ns_0_i_0_0_0_cascade_ ;
    wire \uart_tx.N_187_1_i ;
    wire \uart_tx.M_ctr_qZ0Z_0 ;
    wire bfn_21_4_0_;
    wire \uart_tx.M_ctr_qZ0Z_1 ;
    wire \uart_tx.un1_M_ctr_q_3_cry_0 ;
    wire \uart_tx.un1_M_ctr_q_3_cry_1 ;
    wire \uart_tx.M_ctr_qZ0Z_3 ;
    wire \uart_tx.un1_M_ctr_q_3_cry_2 ;
    wire \uart_tx.M_ctr_qZ0Z_4 ;
    wire \uart_tx.un1_M_ctr_q_3_cry_3 ;
    wire \uart_tx.un1_M_ctr_q_3_cry_4 ;
    wire \uart_tx.un1_M_ctr_q_3_cry_5 ;
    wire \uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_ ;
    wire \uart_tx.M_ctr_qZ0Z_6 ;
    wire usb_tx_c;
    wire \uart_tx.M_txReg_d_0_iv_0_1 ;
    wire \uart_rx.un1_M_ctr_q_5_ac0_1_out ;
    wire \uart_rx.M_bitCtr_q_RNI578A4Z0Z_0_cascade_ ;
    wire \uart_rx.M_ctr_qZ0Z_3 ;
    wire \uart_rx.M_ctr_qZ0Z_5 ;
    wire \uart_rx.M_ctr_qZ0Z_2 ;
    wire \uart_rx.M_ctr_qZ0Z_1 ;
    wire \uart_rx.M_ctr_q_RNIBJBV1Z0Z_1 ;
    wire \uart_rx.M_ctr_qZ0Z_6 ;
    wire \uart_rx.M_ctr_qZ0Z_4 ;
    wire \uart_rx.M_ctr_q_RNIBJBV1Z0Z_1_cascade_ ;
    wire \uart_rx.M_ctr_qZ0Z_0 ;
    wire \uart_rx.M_ctr_q_RNILBSE3Z0Z_6_cascade_ ;
    wire \uart_rx.M_state_q_RNIRDQO7_0Z0Z_0 ;
    wire uart_tx_N_187_1_cascade_;
    wire \uart_tx.N_58 ;
    wire \uart_tx.M_savedData_qZ0Z_0 ;
    wire \uart_tx.M_txReg_d_3_3_i_m4_ns_1_cascade_ ;
    wire \uart_tx.N_66 ;
    wire \uart_tx.M_state_qZ0Z_0 ;
    wire \uart_tx.SUM_i_i_o4_1_1 ;
    wire \uart_tx.SUM_i_i_o4_1_1_cascade_ ;
    wire \uart_tx.M_bitCtr_qZ0Z_0 ;
    wire \uart_tx.M_state_qZ0Z_1 ;
    wire \uart_tx.M_savedData_qZ0Z_3 ;
    wire \uart_tx.M_txReg_d_0_iv_0_a2_1_1_cascade_ ;
    wire \uart_tx.M_bitCtr_qZ0Z_1 ;
    wire \uart_tx.N_81 ;
    wire \uart_tx.M_ctr_q_RNO_0Z0Z_2 ;
    wire \uart_tx.M_ctr_qZ0Z_2 ;
    wire \uart_tx.N_183_0 ;
    wire \uart_tx.N_52_i ;
    wire \uart_tx.M_ctr_q_RNO_0Z0Z_5 ;
    wire \uart_tx.M_ctr_qZ0Z_5 ;
    wire \greeter.M_state_d_0_sqmuxa_1_5_cascade_ ;
    wire \uart_rx.M_state_q_ns_1_cascade_ ;
    wire \uart_rx.M_bitCtr_qZ0Z_2 ;
    wire \uart_rx.M_state_q_37_d ;
    wire \uart_rx.M_state_q_37_d_cascade_ ;
    wire \uart_rx.M_bitCtr_q_RNI578A4Z0Z_0 ;
    wire \uart_rx.M_bitCtr_qZ0Z_1 ;
    wire \uart_rx.M_ctr_q_RNILBSE3Z0Z_6 ;
    wire \uart_rx.M_bitCtr_qZ0Z_0 ;
    wire \greeter.M_state_q_0_cascade_ ;
    wire \greeter.M_state_d_0_sqmuxa_1_7 ;
    wire M_uart_rx_new_data_0;
    wire \greeter.M_state_d_0_sqmuxa_1_6 ;
    wire \uart_tx.M_bitCtr_qZ0Z_2 ;
    wire \uart_tx.N_65 ;
    wire \uart_rx.M_state_qZ0Z_1 ;
    wire \uart_rx.m19_0_o2 ;
    wire M_reset_cond_out_0;
    wire \uart_rx.m19_0_0_cascade_ ;
    wire \uart_rx.M_state_d_0_sqmuxa_1 ;
    wire \uart_rx.M_state_qZ0Z_0 ;
    wire M_greeter_tx_data_0;
    wire N_35_cascade_;
    wire \uart_tx.M_savedData_qZ0Z_6 ;
    wire N_41_cascade_;
    wire \uart_tx.M_savedData_qZ0Z_2 ;
    wire bfn_23_4_0_;
    wire \greeter.un1_M_count_q_1_cry_0 ;
    wire \greeter.un1_M_count_q_1_cry_1 ;
    wire \greeter.un1_M_count_q_1_cry_2 ;
    wire m14_0;
    wire M_greeter_tx_data_4_cascade_;
    wire \uart_tx.M_savedData_qZ0Z_4 ;
    wire M_uart_rx_data_7;
    wire M_uart_rx_data_6;
    wire M_uart_rx_data_0;
    wire M_uart_rx_data_2;
    wire M_uart_rx_data_1;
    wire M_uart_rx_data_5;
    wire M_uart_rx_data_4;
    wire M_uart_rx_data_3;
    wire \uart_rx.N_25_i ;
    wire N_37_cascade_;
    wire \uart_tx.M_savedData_qZ0Z_5 ;
    wire greeter_M_state_q;
    wire M_greeter_tx_data_1_cascade_;
    wire uart_tx_N_187_1;
    wire \uart_tx.M_savedData_qZ1Z_1 ;
    wire \greeter.M_count_qZ1Z_2 ;
    wire \greeter.M_count_qZ0Z_1 ;
    wire \greeter.M_count_qZ0Z_3 ;
    wire \greeter.M_count_qZ0Z_0 ;
    wire \greeter.un1_M_state_d_0_sqmuxa_1_0_a2_0_0 ;
    wire usb_rx_c;
    wire \uart_rx.M_rxd_qZ0 ;
    wire clk_c_g;
    wire _gnd_net_;

    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__3163),
            .GLOBALBUFFEROUTPUT(clk_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__3165),
            .DIN(N__3164),
            .DOUT(N__3163),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__3165),
            .PADOUT(N__3164),
            .PADIN(N__3163),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_0_iopad (
            .OE(N__3154),
            .DIN(N__3153),
            .DOUT(N__3152),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__3154),
            .PADOUT(N__3153),
            .PADIN(N__3152),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_1_iopad (
            .OE(N__3145),
            .DIN(N__3144),
            .DOUT(N__3143),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__3145),
            .PADOUT(N__3144),
            .PADIN(N__3143),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_2_iopad (
            .OE(N__3136),
            .DIN(N__3135),
            .DOUT(N__3134),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__3136),
            .PADOUT(N__3135),
            .PADIN(N__3134),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_3_iopad (
            .OE(N__3127),
            .DIN(N__3126),
            .DOUT(N__3125),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__3127),
            .PADOUT(N__3126),
            .PADIN(N__3125),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_4_iopad (
            .OE(N__3118),
            .DIN(N__3117),
            .DOUT(N__3116),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__3118),
            .PADOUT(N__3117),
            .PADIN(N__3116),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_5_iopad (
            .OE(N__3109),
            .DIN(N__3108),
            .DOUT(N__3107),
            .PACKAGEPIN(led[5]));
    defparam led_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_5_preio (
            .PADOEN(N__3109),
            .PADOUT(N__3108),
            .PADIN(N__3107),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_6_iopad (
            .OE(N__3100),
            .DIN(N__3099),
            .DOUT(N__3098),
            .PACKAGEPIN(led[6]));
    defparam led_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_6_preio (
            .PADOEN(N__3100),
            .PADOUT(N__3099),
            .PADIN(N__3098),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_7_iopad (
            .OE(N__3091),
            .DIN(N__3090),
            .DOUT(N__3089),
            .PACKAGEPIN(led[7]));
    defparam led_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_7_preio (
            .PADOEN(N__3091),
            .PADOUT(N__3090),
            .PADIN(N__3089),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__3082),
            .DIN(N__3081),
            .DOUT(N__3080),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__3082),
            .PADOUT(N__3081),
            .PADIN(N__3080),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD usb_rx_ibuf_iopad (
            .OE(N__3073),
            .DIN(N__3072),
            .DOUT(N__3071),
            .PACKAGEPIN(usb_rx));
    defparam usb_rx_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam usb_rx_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO usb_rx_ibuf_preio (
            .PADOEN(N__3073),
            .PADOUT(N__3072),
            .PADIN(N__3071),
            .CLOCKENABLE(),
            .DIN0(usb_rx_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD usb_tx_obuf_iopad (
            .OE(N__3064),
            .DIN(N__3063),
            .DOUT(N__3062),
            .PACKAGEPIN(usb_tx));
    defparam usb_tx_obuf_preio.NEG_TRIGGER=1'b0;
    defparam usb_tx_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO usb_tx_obuf_preio (
            .PADOEN(N__3064),
            .PADOUT(N__3063),
            .PADIN(N__3062),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__1464),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__694 (
            .O(N__3045),
            .I(N__3041));
    InMux I__693 (
            .O(N__3044),
            .I(N__3038));
    LocalMux I__692 (
            .O(N__3041),
            .I(M_uart_rx_data_4));
    LocalMux I__691 (
            .O(N__3038),
            .I(M_uart_rx_data_4));
    InMux I__690 (
            .O(N__3033),
            .I(N__3029));
    InMux I__689 (
            .O(N__3032),
            .I(N__3026));
    LocalMux I__688 (
            .O(N__3029),
            .I(M_uart_rx_data_3));
    LocalMux I__687 (
            .O(N__3026),
            .I(M_uart_rx_data_3));
    CEMux I__686 (
            .O(N__3021),
            .I(N__3018));
    LocalMux I__685 (
            .O(N__3018),
            .I(N__3014));
    CEMux I__684 (
            .O(N__3017),
            .I(N__3011));
    Span4Mux_v I__683 (
            .O(N__3014),
            .I(N__3006));
    LocalMux I__682 (
            .O(N__3011),
            .I(N__3006));
    Span4Mux_s0_v I__681 (
            .O(N__3006),
            .I(N__3003));
    Odrv4 I__680 (
            .O(N__3003),
            .I(\uart_rx.N_25_i ));
    CascadeMux I__679 (
            .O(N__3000),
            .I(N_37_cascade_));
    InMux I__678 (
            .O(N__2997),
            .I(N__2993));
    InMux I__677 (
            .O(N__2996),
            .I(N__2990));
    LocalMux I__676 (
            .O(N__2993),
            .I(\uart_tx.M_savedData_qZ0Z_5 ));
    LocalMux I__675 (
            .O(N__2990),
            .I(\uart_tx.M_savedData_qZ0Z_5 ));
    CascadeMux I__674 (
            .O(N__2985),
            .I(N__2981));
    CascadeMux I__673 (
            .O(N__2984),
            .I(N__2978));
    InMux I__672 (
            .O(N__2981),
            .I(N__2969));
    InMux I__671 (
            .O(N__2978),
            .I(N__2966));
    CascadeMux I__670 (
            .O(N__2977),
            .I(N__2961));
    InMux I__669 (
            .O(N__2976),
            .I(N__2954));
    InMux I__668 (
            .O(N__2975),
            .I(N__2954));
    InMux I__667 (
            .O(N__2974),
            .I(N__2947));
    InMux I__666 (
            .O(N__2973),
            .I(N__2947));
    InMux I__665 (
            .O(N__2972),
            .I(N__2947));
    LocalMux I__664 (
            .O(N__2969),
            .I(N__2944));
    LocalMux I__663 (
            .O(N__2966),
            .I(N__2941));
    InMux I__662 (
            .O(N__2965),
            .I(N__2934));
    InMux I__661 (
            .O(N__2964),
            .I(N__2934));
    InMux I__660 (
            .O(N__2961),
            .I(N__2931));
    InMux I__659 (
            .O(N__2960),
            .I(N__2926));
    InMux I__658 (
            .O(N__2959),
            .I(N__2926));
    LocalMux I__657 (
            .O(N__2954),
            .I(N__2921));
    LocalMux I__656 (
            .O(N__2947),
            .I(N__2921));
    Span4Mux_v I__655 (
            .O(N__2944),
            .I(N__2916));
    Span4Mux_h I__654 (
            .O(N__2941),
            .I(N__2916));
    InMux I__653 (
            .O(N__2940),
            .I(N__2913));
    InMux I__652 (
            .O(N__2939),
            .I(N__2910));
    LocalMux I__651 (
            .O(N__2934),
            .I(greeter_M_state_q));
    LocalMux I__650 (
            .O(N__2931),
            .I(greeter_M_state_q));
    LocalMux I__649 (
            .O(N__2926),
            .I(greeter_M_state_q));
    Odrv4 I__648 (
            .O(N__2921),
            .I(greeter_M_state_q));
    Odrv4 I__647 (
            .O(N__2916),
            .I(greeter_M_state_q));
    LocalMux I__646 (
            .O(N__2913),
            .I(greeter_M_state_q));
    LocalMux I__645 (
            .O(N__2910),
            .I(greeter_M_state_q));
    CascadeMux I__644 (
            .O(N__2895),
            .I(M_greeter_tx_data_1_cascade_));
    SRMux I__643 (
            .O(N__2892),
            .I(N__2889));
    LocalMux I__642 (
            .O(N__2889),
            .I(N__2881));
    InMux I__641 (
            .O(N__2888),
            .I(N__2865));
    InMux I__640 (
            .O(N__2887),
            .I(N__2865));
    InMux I__639 (
            .O(N__2886),
            .I(N__2860));
    InMux I__638 (
            .O(N__2885),
            .I(N__2860));
    CascadeMux I__637 (
            .O(N__2884),
            .I(N__2855));
    Span4Mux_h I__636 (
            .O(N__2881),
            .I(N__2852));
    InMux I__635 (
            .O(N__2880),
            .I(N__2849));
    InMux I__634 (
            .O(N__2879),
            .I(N__2842));
    InMux I__633 (
            .O(N__2878),
            .I(N__2842));
    InMux I__632 (
            .O(N__2877),
            .I(N__2842));
    InMux I__631 (
            .O(N__2876),
            .I(N__2837));
    InMux I__630 (
            .O(N__2875),
            .I(N__2837));
    InMux I__629 (
            .O(N__2874),
            .I(N__2832));
    InMux I__628 (
            .O(N__2873),
            .I(N__2832));
    InMux I__627 (
            .O(N__2872),
            .I(N__2825));
    InMux I__626 (
            .O(N__2871),
            .I(N__2825));
    InMux I__625 (
            .O(N__2870),
            .I(N__2825));
    LocalMux I__624 (
            .O(N__2865),
            .I(N__2820));
    LocalMux I__623 (
            .O(N__2860),
            .I(N__2820));
    InMux I__622 (
            .O(N__2859),
            .I(N__2817));
    InMux I__621 (
            .O(N__2858),
            .I(N__2812));
    InMux I__620 (
            .O(N__2855),
            .I(N__2812));
    Span4Mux_s0_v I__619 (
            .O(N__2852),
            .I(N__2809));
    LocalMux I__618 (
            .O(N__2849),
            .I(uart_tx_N_187_1));
    LocalMux I__617 (
            .O(N__2842),
            .I(uart_tx_N_187_1));
    LocalMux I__616 (
            .O(N__2837),
            .I(uart_tx_N_187_1));
    LocalMux I__615 (
            .O(N__2832),
            .I(uart_tx_N_187_1));
    LocalMux I__614 (
            .O(N__2825),
            .I(uart_tx_N_187_1));
    Odrv4 I__613 (
            .O(N__2820),
            .I(uart_tx_N_187_1));
    LocalMux I__612 (
            .O(N__2817),
            .I(uart_tx_N_187_1));
    LocalMux I__611 (
            .O(N__2812),
            .I(uart_tx_N_187_1));
    Odrv4 I__610 (
            .O(N__2809),
            .I(uart_tx_N_187_1));
    InMux I__609 (
            .O(N__2790),
            .I(N__2786));
    InMux I__608 (
            .O(N__2789),
            .I(N__2783));
    LocalMux I__607 (
            .O(N__2786),
            .I(\uart_tx.M_savedData_qZ1Z_1 ));
    LocalMux I__606 (
            .O(N__2783),
            .I(\uart_tx.M_savedData_qZ1Z_1 ));
    CascadeMux I__605 (
            .O(N__2778),
            .I(N__2768));
    CascadeMux I__604 (
            .O(N__2777),
            .I(N__2765));
    InMux I__603 (
            .O(N__2776),
            .I(N__2757));
    InMux I__602 (
            .O(N__2775),
            .I(N__2757));
    InMux I__601 (
            .O(N__2774),
            .I(N__2757));
    InMux I__600 (
            .O(N__2773),
            .I(N__2750));
    InMux I__599 (
            .O(N__2772),
            .I(N__2750));
    InMux I__598 (
            .O(N__2771),
            .I(N__2750));
    InMux I__597 (
            .O(N__2768),
            .I(N__2743));
    InMux I__596 (
            .O(N__2765),
            .I(N__2743));
    InMux I__595 (
            .O(N__2764),
            .I(N__2743));
    LocalMux I__594 (
            .O(N__2757),
            .I(N__2740));
    LocalMux I__593 (
            .O(N__2750),
            .I(\greeter.M_count_qZ1Z_2 ));
    LocalMux I__592 (
            .O(N__2743),
            .I(\greeter.M_count_qZ1Z_2 ));
    Odrv4 I__591 (
            .O(N__2740),
            .I(\greeter.M_count_qZ1Z_2 ));
    CascadeMux I__590 (
            .O(N__2733),
            .I(N__2729));
    InMux I__589 (
            .O(N__2732),
            .I(N__2715));
    InMux I__588 (
            .O(N__2729),
            .I(N__2715));
    InMux I__587 (
            .O(N__2728),
            .I(N__2715));
    InMux I__586 (
            .O(N__2727),
            .I(N__2708));
    InMux I__585 (
            .O(N__2726),
            .I(N__2708));
    InMux I__584 (
            .O(N__2725),
            .I(N__2708));
    InMux I__583 (
            .O(N__2724),
            .I(N__2701));
    InMux I__582 (
            .O(N__2723),
            .I(N__2701));
    InMux I__581 (
            .O(N__2722),
            .I(N__2701));
    LocalMux I__580 (
            .O(N__2715),
            .I(\greeter.M_count_qZ0Z_1 ));
    LocalMux I__579 (
            .O(N__2708),
            .I(\greeter.M_count_qZ0Z_1 ));
    LocalMux I__578 (
            .O(N__2701),
            .I(\greeter.M_count_qZ0Z_1 ));
    CascadeMux I__577 (
            .O(N__2694),
            .I(N__2686));
    CascadeMux I__576 (
            .O(N__2693),
            .I(N__2680));
    CascadeMux I__575 (
            .O(N__2692),
            .I(N__2677));
    CascadeMux I__574 (
            .O(N__2691),
            .I(N__2674));
    CascadeMux I__573 (
            .O(N__2690),
            .I(N__2671));
    InMux I__572 (
            .O(N__2689),
            .I(N__2664));
    InMux I__571 (
            .O(N__2686),
            .I(N__2664));
    InMux I__570 (
            .O(N__2685),
            .I(N__2664));
    InMux I__569 (
            .O(N__2684),
            .I(N__2657));
    InMux I__568 (
            .O(N__2683),
            .I(N__2657));
    InMux I__567 (
            .O(N__2680),
            .I(N__2657));
    InMux I__566 (
            .O(N__2677),
            .I(N__2650));
    InMux I__565 (
            .O(N__2674),
            .I(N__2650));
    InMux I__564 (
            .O(N__2671),
            .I(N__2650));
    LocalMux I__563 (
            .O(N__2664),
            .I(\greeter.M_count_qZ0Z_3 ));
    LocalMux I__562 (
            .O(N__2657),
            .I(\greeter.M_count_qZ0Z_3 ));
    LocalMux I__561 (
            .O(N__2650),
            .I(\greeter.M_count_qZ0Z_3 ));
    InMux I__560 (
            .O(N__2643),
            .I(N__2632));
    InMux I__559 (
            .O(N__2642),
            .I(N__2627));
    InMux I__558 (
            .O(N__2641),
            .I(N__2627));
    InMux I__557 (
            .O(N__2640),
            .I(N__2620));
    InMux I__556 (
            .O(N__2639),
            .I(N__2620));
    InMux I__555 (
            .O(N__2638),
            .I(N__2620));
    InMux I__554 (
            .O(N__2637),
            .I(N__2613));
    InMux I__553 (
            .O(N__2636),
            .I(N__2613));
    InMux I__552 (
            .O(N__2635),
            .I(N__2613));
    LocalMux I__551 (
            .O(N__2632),
            .I(\greeter.M_count_qZ0Z_0 ));
    LocalMux I__550 (
            .O(N__2627),
            .I(\greeter.M_count_qZ0Z_0 ));
    LocalMux I__549 (
            .O(N__2620),
            .I(\greeter.M_count_qZ0Z_0 ));
    LocalMux I__548 (
            .O(N__2613),
            .I(\greeter.M_count_qZ0Z_0 ));
    InMux I__547 (
            .O(N__2604),
            .I(N__2601));
    LocalMux I__546 (
            .O(N__2601),
            .I(\greeter.un1_M_state_d_0_sqmuxa_1_0_a2_0_0 ));
    InMux I__545 (
            .O(N__2598),
            .I(N__2595));
    LocalMux I__544 (
            .O(N__2595),
            .I(N__2592));
    Odrv12 I__543 (
            .O(N__2592),
            .I(usb_rx_c));
    CascadeMux I__542 (
            .O(N__2589),
            .I(N__2585));
    InMux I__541 (
            .O(N__2588),
            .I(N__2581));
    InMux I__540 (
            .O(N__2585),
            .I(N__2578));
    CascadeMux I__539 (
            .O(N__2584),
            .I(N__2575));
    LocalMux I__538 (
            .O(N__2581),
            .I(N__2572));
    LocalMux I__537 (
            .O(N__2578),
            .I(N__2569));
    InMux I__536 (
            .O(N__2575),
            .I(N__2566));
    Span4Mux_h I__535 (
            .O(N__2572),
            .I(N__2563));
    Span4Mux_v I__534 (
            .O(N__2569),
            .I(N__2558));
    LocalMux I__533 (
            .O(N__2566),
            .I(N__2558));
    Odrv4 I__532 (
            .O(N__2563),
            .I(\uart_rx.M_rxd_qZ0 ));
    Odrv4 I__531 (
            .O(N__2558),
            .I(\uart_rx.M_rxd_qZ0 ));
    ClkMux I__530 (
            .O(N__2553),
            .I(N__2508));
    ClkMux I__529 (
            .O(N__2552),
            .I(N__2508));
    ClkMux I__528 (
            .O(N__2551),
            .I(N__2508));
    ClkMux I__527 (
            .O(N__2550),
            .I(N__2508));
    ClkMux I__526 (
            .O(N__2549),
            .I(N__2508));
    ClkMux I__525 (
            .O(N__2548),
            .I(N__2508));
    ClkMux I__524 (
            .O(N__2547),
            .I(N__2508));
    ClkMux I__523 (
            .O(N__2546),
            .I(N__2508));
    ClkMux I__522 (
            .O(N__2545),
            .I(N__2508));
    ClkMux I__521 (
            .O(N__2544),
            .I(N__2508));
    ClkMux I__520 (
            .O(N__2543),
            .I(N__2508));
    ClkMux I__519 (
            .O(N__2542),
            .I(N__2508));
    ClkMux I__518 (
            .O(N__2541),
            .I(N__2508));
    ClkMux I__517 (
            .O(N__2540),
            .I(N__2508));
    ClkMux I__516 (
            .O(N__2539),
            .I(N__2508));
    GlobalMux I__515 (
            .O(N__2508),
            .I(N__2505));
    gio2CtrlBuf I__514 (
            .O(N__2505),
            .I(clk_c_g));
    CascadeMux I__513 (
            .O(N__2502),
            .I(M_greeter_tx_data_4_cascade_));
    CascadeMux I__512 (
            .O(N__2499),
            .I(N__2495));
    InMux I__511 (
            .O(N__2498),
            .I(N__2492));
    InMux I__510 (
            .O(N__2495),
            .I(N__2489));
    LocalMux I__509 (
            .O(N__2492),
            .I(\uart_tx.M_savedData_qZ0Z_4 ));
    LocalMux I__508 (
            .O(N__2489),
            .I(\uart_tx.M_savedData_qZ0Z_4 ));
    CascadeMux I__507 (
            .O(N__2484),
            .I(N__2480));
    InMux I__506 (
            .O(N__2483),
            .I(N__2477));
    InMux I__505 (
            .O(N__2480),
            .I(N__2474));
    LocalMux I__504 (
            .O(N__2477),
            .I(M_uart_rx_data_7));
    LocalMux I__503 (
            .O(N__2474),
            .I(M_uart_rx_data_7));
    InMux I__502 (
            .O(N__2469),
            .I(N__2465));
    InMux I__501 (
            .O(N__2468),
            .I(N__2462));
    LocalMux I__500 (
            .O(N__2465),
            .I(M_uart_rx_data_6));
    LocalMux I__499 (
            .O(N__2462),
            .I(M_uart_rx_data_6));
    InMux I__498 (
            .O(N__2457),
            .I(N__2454));
    LocalMux I__497 (
            .O(N__2454),
            .I(M_uart_rx_data_0));
    InMux I__496 (
            .O(N__2451),
            .I(N__2447));
    InMux I__495 (
            .O(N__2450),
            .I(N__2444));
    LocalMux I__494 (
            .O(N__2447),
            .I(M_uart_rx_data_2));
    LocalMux I__493 (
            .O(N__2444),
            .I(M_uart_rx_data_2));
    InMux I__492 (
            .O(N__2439),
            .I(N__2435));
    InMux I__491 (
            .O(N__2438),
            .I(N__2432));
    LocalMux I__490 (
            .O(N__2435),
            .I(M_uart_rx_data_1));
    LocalMux I__489 (
            .O(N__2432),
            .I(M_uart_rx_data_1));
    InMux I__488 (
            .O(N__2427),
            .I(N__2423));
    InMux I__487 (
            .O(N__2426),
            .I(N__2420));
    LocalMux I__486 (
            .O(N__2423),
            .I(M_uart_rx_data_5));
    LocalMux I__485 (
            .O(N__2420),
            .I(M_uart_rx_data_5));
    CascadeMux I__484 (
            .O(N__2415),
            .I(N_35_cascade_));
    InMux I__483 (
            .O(N__2412),
            .I(N__2408));
    InMux I__482 (
            .O(N__2411),
            .I(N__2405));
    LocalMux I__481 (
            .O(N__2408),
            .I(\uart_tx.M_savedData_qZ0Z_6 ));
    LocalMux I__480 (
            .O(N__2405),
            .I(\uart_tx.M_savedData_qZ0Z_6 ));
    CascadeMux I__479 (
            .O(N__2400),
            .I(N_41_cascade_));
    InMux I__478 (
            .O(N__2397),
            .I(N__2393));
    InMux I__477 (
            .O(N__2396),
            .I(N__2390));
    LocalMux I__476 (
            .O(N__2393),
            .I(N__2385));
    LocalMux I__475 (
            .O(N__2390),
            .I(N__2385));
    Odrv4 I__474 (
            .O(N__2385),
            .I(\uart_tx.M_savedData_qZ0Z_2 ));
    InMux I__473 (
            .O(N__2382),
            .I(\greeter.un1_M_count_q_1_cry_0 ));
    InMux I__472 (
            .O(N__2379),
            .I(\greeter.un1_M_count_q_1_cry_1 ));
    InMux I__471 (
            .O(N__2376),
            .I(\greeter.un1_M_count_q_1_cry_2 ));
    InMux I__470 (
            .O(N__2373),
            .I(N__2370));
    LocalMux I__469 (
            .O(N__2370),
            .I(m14_0));
    CascadeMux I__468 (
            .O(N__2367),
            .I(\uart_rx.M_state_q_37_d_cascade_ ));
    InMux I__467 (
            .O(N__2364),
            .I(N__2355));
    InMux I__466 (
            .O(N__2363),
            .I(N__2355));
    InMux I__465 (
            .O(N__2362),
            .I(N__2355));
    LocalMux I__464 (
            .O(N__2355),
            .I(\uart_rx.M_bitCtr_q_RNI578A4Z0Z_0 ));
    CascadeMux I__463 (
            .O(N__2352),
            .I(N__2348));
    InMux I__462 (
            .O(N__2351),
            .I(N__2339));
    InMux I__461 (
            .O(N__2348),
            .I(N__2339));
    InMux I__460 (
            .O(N__2347),
            .I(N__2339));
    InMux I__459 (
            .O(N__2346),
            .I(N__2336));
    LocalMux I__458 (
            .O(N__2339),
            .I(\uart_rx.M_bitCtr_qZ0Z_1 ));
    LocalMux I__457 (
            .O(N__2336),
            .I(\uart_rx.M_bitCtr_qZ0Z_1 ));
    InMux I__456 (
            .O(N__2331),
            .I(N__2325));
    InMux I__455 (
            .O(N__2330),
            .I(N__2322));
    InMux I__454 (
            .O(N__2329),
            .I(N__2319));
    InMux I__453 (
            .O(N__2328),
            .I(N__2316));
    LocalMux I__452 (
            .O(N__2325),
            .I(\uart_rx.M_ctr_q_RNILBSE3Z0Z_6 ));
    LocalMux I__451 (
            .O(N__2322),
            .I(\uart_rx.M_ctr_q_RNILBSE3Z0Z_6 ));
    LocalMux I__450 (
            .O(N__2319),
            .I(\uart_rx.M_ctr_q_RNILBSE3Z0Z_6 ));
    LocalMux I__449 (
            .O(N__2316),
            .I(\uart_rx.M_ctr_q_RNILBSE3Z0Z_6 ));
    InMux I__448 (
            .O(N__2307),
            .I(N__2303));
    InMux I__447 (
            .O(N__2306),
            .I(N__2300));
    LocalMux I__446 (
            .O(N__2303),
            .I(\uart_rx.M_bitCtr_qZ0Z_0 ));
    LocalMux I__445 (
            .O(N__2300),
            .I(\uart_rx.M_bitCtr_qZ0Z_0 ));
    CascadeMux I__444 (
            .O(N__2295),
            .I(\greeter.M_state_q_0_cascade_ ));
    InMux I__443 (
            .O(N__2292),
            .I(N__2289));
    LocalMux I__442 (
            .O(N__2289),
            .I(N__2286));
    Odrv4 I__441 (
            .O(N__2286),
            .I(\greeter.M_state_d_0_sqmuxa_1_7 ));
    CascadeMux I__440 (
            .O(N__2283),
            .I(N__2280));
    InMux I__439 (
            .O(N__2280),
            .I(N__2277));
    LocalMux I__438 (
            .O(N__2277),
            .I(M_uart_rx_new_data_0));
    InMux I__437 (
            .O(N__2274),
            .I(N__2271));
    LocalMux I__436 (
            .O(N__2271),
            .I(\greeter.M_state_d_0_sqmuxa_1_6 ));
    InMux I__435 (
            .O(N__2268),
            .I(N__2261));
    InMux I__434 (
            .O(N__2267),
            .I(N__2258));
    InMux I__433 (
            .O(N__2266),
            .I(N__2255));
    InMux I__432 (
            .O(N__2265),
            .I(N__2250));
    InMux I__431 (
            .O(N__2264),
            .I(N__2250));
    LocalMux I__430 (
            .O(N__2261),
            .I(\uart_tx.M_bitCtr_qZ0Z_2 ));
    LocalMux I__429 (
            .O(N__2258),
            .I(\uart_tx.M_bitCtr_qZ0Z_2 ));
    LocalMux I__428 (
            .O(N__2255),
            .I(\uart_tx.M_bitCtr_qZ0Z_2 ));
    LocalMux I__427 (
            .O(N__2250),
            .I(\uart_tx.M_bitCtr_qZ0Z_2 ));
    CascadeMux I__426 (
            .O(N__2241),
            .I(N__2238));
    InMux I__425 (
            .O(N__2238),
            .I(N__2235));
    LocalMux I__424 (
            .O(N__2235),
            .I(\uart_tx.N_65 ));
    CascadeMux I__423 (
            .O(N__2232),
            .I(N__2229));
    InMux I__422 (
            .O(N__2229),
            .I(N__2223));
    CascadeMux I__421 (
            .O(N__2228),
            .I(N__2220));
    InMux I__420 (
            .O(N__2227),
            .I(N__2217));
    CascadeMux I__419 (
            .O(N__2226),
            .I(N__2213));
    LocalMux I__418 (
            .O(N__2223),
            .I(N__2209));
    InMux I__417 (
            .O(N__2220),
            .I(N__2204));
    LocalMux I__416 (
            .O(N__2217),
            .I(N__2201));
    InMux I__415 (
            .O(N__2216),
            .I(N__2198));
    InMux I__414 (
            .O(N__2213),
            .I(N__2193));
    InMux I__413 (
            .O(N__2212),
            .I(N__2193));
    Span4Mux_v I__412 (
            .O(N__2209),
            .I(N__2190));
    InMux I__411 (
            .O(N__2208),
            .I(N__2185));
    InMux I__410 (
            .O(N__2207),
            .I(N__2185));
    LocalMux I__409 (
            .O(N__2204),
            .I(\uart_rx.M_state_qZ0Z_1 ));
    Odrv12 I__408 (
            .O(N__2201),
            .I(\uart_rx.M_state_qZ0Z_1 ));
    LocalMux I__407 (
            .O(N__2198),
            .I(\uart_rx.M_state_qZ0Z_1 ));
    LocalMux I__406 (
            .O(N__2193),
            .I(\uart_rx.M_state_qZ0Z_1 ));
    Odrv4 I__405 (
            .O(N__2190),
            .I(\uart_rx.M_state_qZ0Z_1 ));
    LocalMux I__404 (
            .O(N__2185),
            .I(\uart_rx.M_state_qZ0Z_1 ));
    InMux I__403 (
            .O(N__2172),
            .I(N__2166));
    InMux I__402 (
            .O(N__2171),
            .I(N__2163));
    InMux I__401 (
            .O(N__2170),
            .I(N__2160));
    InMux I__400 (
            .O(N__2169),
            .I(N__2157));
    LocalMux I__399 (
            .O(N__2166),
            .I(\uart_rx.m19_0_o2 ));
    LocalMux I__398 (
            .O(N__2163),
            .I(\uart_rx.m19_0_o2 ));
    LocalMux I__397 (
            .O(N__2160),
            .I(\uart_rx.m19_0_o2 ));
    LocalMux I__396 (
            .O(N__2157),
            .I(\uart_rx.m19_0_o2 ));
    InMux I__395 (
            .O(N__2148),
            .I(N__2144));
    InMux I__394 (
            .O(N__2147),
            .I(N__2141));
    LocalMux I__393 (
            .O(N__2144),
            .I(N__2135));
    LocalMux I__392 (
            .O(N__2141),
            .I(N__2132));
    InMux I__391 (
            .O(N__2140),
            .I(N__2129));
    InMux I__390 (
            .O(N__2139),
            .I(N__2124));
    InMux I__389 (
            .O(N__2138),
            .I(N__2124));
    Span4Mux_s1_v I__388 (
            .O(N__2135),
            .I(N__2117));
    Span4Mux_v I__387 (
            .O(N__2132),
            .I(N__2117));
    LocalMux I__386 (
            .O(N__2129),
            .I(N__2117));
    LocalMux I__385 (
            .O(N__2124),
            .I(N__2114));
    Odrv4 I__384 (
            .O(N__2117),
            .I(M_reset_cond_out_0));
    Odrv4 I__383 (
            .O(N__2114),
            .I(M_reset_cond_out_0));
    CascadeMux I__382 (
            .O(N__2109),
            .I(\uart_rx.m19_0_0_cascade_ ));
    InMux I__381 (
            .O(N__2106),
            .I(N__2103));
    LocalMux I__380 (
            .O(N__2103),
            .I(\uart_rx.M_state_d_0_sqmuxa_1 ));
    InMux I__379 (
            .O(N__2100),
            .I(N__2096));
    InMux I__378 (
            .O(N__2099),
            .I(N__2087));
    LocalMux I__377 (
            .O(N__2096),
            .I(N__2084));
    InMux I__376 (
            .O(N__2095),
            .I(N__2081));
    InMux I__375 (
            .O(N__2094),
            .I(N__2076));
    InMux I__374 (
            .O(N__2093),
            .I(N__2076));
    InMux I__373 (
            .O(N__2092),
            .I(N__2073));
    InMux I__372 (
            .O(N__2091),
            .I(N__2070));
    InMux I__371 (
            .O(N__2090),
            .I(N__2067));
    LocalMux I__370 (
            .O(N__2087),
            .I(N__2062));
    Span4Mux_s2_v I__369 (
            .O(N__2084),
            .I(N__2062));
    LocalMux I__368 (
            .O(N__2081),
            .I(N__2057));
    LocalMux I__367 (
            .O(N__2076),
            .I(N__2057));
    LocalMux I__366 (
            .O(N__2073),
            .I(\uart_rx.M_state_qZ0Z_0 ));
    LocalMux I__365 (
            .O(N__2070),
            .I(\uart_rx.M_state_qZ0Z_0 ));
    LocalMux I__364 (
            .O(N__2067),
            .I(\uart_rx.M_state_qZ0Z_0 ));
    Odrv4 I__363 (
            .O(N__2062),
            .I(\uart_rx.M_state_qZ0Z_0 ));
    Odrv4 I__362 (
            .O(N__2057),
            .I(\uart_rx.M_state_qZ0Z_0 ));
    InMux I__361 (
            .O(N__2046),
            .I(N__2043));
    LocalMux I__360 (
            .O(N__2043),
            .I(M_greeter_tx_data_0));
    InMux I__359 (
            .O(N__2040),
            .I(N__2029));
    InMux I__358 (
            .O(N__2039),
            .I(N__2029));
    InMux I__357 (
            .O(N__2038),
            .I(N__2026));
    InMux I__356 (
            .O(N__2037),
            .I(N__2021));
    InMux I__355 (
            .O(N__2036),
            .I(N__2021));
    InMux I__354 (
            .O(N__2035),
            .I(N__2016));
    InMux I__353 (
            .O(N__2034),
            .I(N__2016));
    LocalMux I__352 (
            .O(N__2029),
            .I(\uart_tx.N_183_0 ));
    LocalMux I__351 (
            .O(N__2026),
            .I(\uart_tx.N_183_0 ));
    LocalMux I__350 (
            .O(N__2021),
            .I(\uart_tx.N_183_0 ));
    LocalMux I__349 (
            .O(N__2016),
            .I(\uart_tx.N_183_0 ));
    CascadeMux I__348 (
            .O(N__2007),
            .I(N__2004));
    InMux I__347 (
            .O(N__2004),
            .I(N__1999));
    CascadeMux I__346 (
            .O(N__2003),
            .I(N__1995));
    CascadeMux I__345 (
            .O(N__2002),
            .I(N__1992));
    LocalMux I__344 (
            .O(N__1999),
            .I(N__1989));
    InMux I__343 (
            .O(N__1998),
            .I(N__1986));
    InMux I__342 (
            .O(N__1995),
            .I(N__1981));
    InMux I__341 (
            .O(N__1992),
            .I(N__1981));
    Span4Mux_h I__340 (
            .O(N__1989),
            .I(N__1976));
    LocalMux I__339 (
            .O(N__1986),
            .I(N__1976));
    LocalMux I__338 (
            .O(N__1981),
            .I(\uart_tx.N_52_i ));
    Odrv4 I__337 (
            .O(N__1976),
            .I(\uart_tx.N_52_i ));
    InMux I__336 (
            .O(N__1971),
            .I(N__1968));
    LocalMux I__335 (
            .O(N__1968),
            .I(\uart_tx.M_ctr_q_RNO_0Z0Z_5 ));
    InMux I__334 (
            .O(N__1965),
            .I(N__1961));
    InMux I__333 (
            .O(N__1964),
            .I(N__1958));
    LocalMux I__332 (
            .O(N__1961),
            .I(N__1955));
    LocalMux I__331 (
            .O(N__1958),
            .I(\uart_tx.M_ctr_qZ0Z_5 ));
    Odrv4 I__330 (
            .O(N__1955),
            .I(\uart_tx.M_ctr_qZ0Z_5 ));
    CascadeMux I__329 (
            .O(N__1950),
            .I(\greeter.M_state_d_0_sqmuxa_1_5_cascade_ ));
    CascadeMux I__328 (
            .O(N__1947),
            .I(\uart_rx.M_state_q_ns_1_cascade_ ));
    InMux I__327 (
            .O(N__1944),
            .I(N__1937));
    InMux I__326 (
            .O(N__1943),
            .I(N__1937));
    InMux I__325 (
            .O(N__1942),
            .I(N__1934));
    LocalMux I__324 (
            .O(N__1937),
            .I(\uart_rx.M_bitCtr_qZ0Z_2 ));
    LocalMux I__323 (
            .O(N__1934),
            .I(\uart_rx.M_bitCtr_qZ0Z_2 ));
    InMux I__322 (
            .O(N__1929),
            .I(N__1926));
    LocalMux I__321 (
            .O(N__1926),
            .I(\uart_rx.M_state_q_37_d ));
    InMux I__320 (
            .O(N__1923),
            .I(N__1917));
    InMux I__319 (
            .O(N__1922),
            .I(N__1917));
    LocalMux I__318 (
            .O(N__1917),
            .I(\uart_tx.M_savedData_qZ0Z_0 ));
    CascadeMux I__317 (
            .O(N__1914),
            .I(\uart_tx.M_txReg_d_3_3_i_m4_ns_1_cascade_ ));
    InMux I__316 (
            .O(N__1911),
            .I(N__1908));
    LocalMux I__315 (
            .O(N__1908),
            .I(\uart_tx.N_66 ));
    CascadeMux I__314 (
            .O(N__1905),
            .I(N__1900));
    CascadeMux I__313 (
            .O(N__1904),
            .I(N__1897));
    CascadeMux I__312 (
            .O(N__1903),
            .I(N__1891));
    InMux I__311 (
            .O(N__1900),
            .I(N__1887));
    InMux I__310 (
            .O(N__1897),
            .I(N__1882));
    InMux I__309 (
            .O(N__1896),
            .I(N__1882));
    InMux I__308 (
            .O(N__1895),
            .I(N__1873));
    InMux I__307 (
            .O(N__1894),
            .I(N__1873));
    InMux I__306 (
            .O(N__1891),
            .I(N__1873));
    InMux I__305 (
            .O(N__1890),
            .I(N__1873));
    LocalMux I__304 (
            .O(N__1887),
            .I(\uart_tx.M_state_qZ0Z_0 ));
    LocalMux I__303 (
            .O(N__1882),
            .I(\uart_tx.M_state_qZ0Z_0 ));
    LocalMux I__302 (
            .O(N__1873),
            .I(\uart_tx.M_state_qZ0Z_0 ));
    InMux I__301 (
            .O(N__1866),
            .I(N__1863));
    LocalMux I__300 (
            .O(N__1863),
            .I(\uart_tx.SUM_i_i_o4_1_1 ));
    CascadeMux I__299 (
            .O(N__1860),
            .I(\uart_tx.SUM_i_i_o4_1_1_cascade_ ));
    InMux I__298 (
            .O(N__1857),
            .I(N__1854));
    LocalMux I__297 (
            .O(N__1854),
            .I(N__1848));
    InMux I__296 (
            .O(N__1853),
            .I(N__1845));
    InMux I__295 (
            .O(N__1852),
            .I(N__1840));
    InMux I__294 (
            .O(N__1851),
            .I(N__1840));
    Odrv4 I__293 (
            .O(N__1848),
            .I(\uart_tx.M_bitCtr_qZ0Z_0 ));
    LocalMux I__292 (
            .O(N__1845),
            .I(\uart_tx.M_bitCtr_qZ0Z_0 ));
    LocalMux I__291 (
            .O(N__1840),
            .I(\uart_tx.M_bitCtr_qZ0Z_0 ));
    CascadeMux I__290 (
            .O(N__1833),
            .I(N__1829));
    InMux I__289 (
            .O(N__1832),
            .I(N__1826));
    InMux I__288 (
            .O(N__1829),
            .I(N__1816));
    LocalMux I__287 (
            .O(N__1826),
            .I(N__1813));
    InMux I__286 (
            .O(N__1825),
            .I(N__1810));
    InMux I__285 (
            .O(N__1824),
            .I(N__1805));
    InMux I__284 (
            .O(N__1823),
            .I(N__1805));
    InMux I__283 (
            .O(N__1822),
            .I(N__1802));
    InMux I__282 (
            .O(N__1821),
            .I(N__1795));
    InMux I__281 (
            .O(N__1820),
            .I(N__1795));
    InMux I__280 (
            .O(N__1819),
            .I(N__1795));
    LocalMux I__279 (
            .O(N__1816),
            .I(\uart_tx.M_state_qZ0Z_1 ));
    Odrv4 I__278 (
            .O(N__1813),
            .I(\uart_tx.M_state_qZ0Z_1 ));
    LocalMux I__277 (
            .O(N__1810),
            .I(\uart_tx.M_state_qZ0Z_1 ));
    LocalMux I__276 (
            .O(N__1805),
            .I(\uart_tx.M_state_qZ0Z_1 ));
    LocalMux I__275 (
            .O(N__1802),
            .I(\uart_tx.M_state_qZ0Z_1 ));
    LocalMux I__274 (
            .O(N__1795),
            .I(\uart_tx.M_state_qZ0Z_1 ));
    InMux I__273 (
            .O(N__1782),
            .I(N__1776));
    InMux I__272 (
            .O(N__1781),
            .I(N__1776));
    LocalMux I__271 (
            .O(N__1776),
            .I(\uart_tx.M_savedData_qZ0Z_3 ));
    CascadeMux I__270 (
            .O(N__1773),
            .I(\uart_tx.M_txReg_d_0_iv_0_a2_1_1_cascade_ ));
    InMux I__269 (
            .O(N__1770),
            .I(N__1767));
    LocalMux I__268 (
            .O(N__1767),
            .I(N__1759));
    InMux I__267 (
            .O(N__1766),
            .I(N__1756));
    InMux I__266 (
            .O(N__1765),
            .I(N__1753));
    InMux I__265 (
            .O(N__1764),
            .I(N__1746));
    InMux I__264 (
            .O(N__1763),
            .I(N__1746));
    InMux I__263 (
            .O(N__1762),
            .I(N__1746));
    Odrv4 I__262 (
            .O(N__1759),
            .I(\uart_tx.M_bitCtr_qZ0Z_1 ));
    LocalMux I__261 (
            .O(N__1756),
            .I(\uart_tx.M_bitCtr_qZ0Z_1 ));
    LocalMux I__260 (
            .O(N__1753),
            .I(\uart_tx.M_bitCtr_qZ0Z_1 ));
    LocalMux I__259 (
            .O(N__1746),
            .I(\uart_tx.M_bitCtr_qZ0Z_1 ));
    InMux I__258 (
            .O(N__1737),
            .I(N__1734));
    LocalMux I__257 (
            .O(N__1734),
            .I(N__1731));
    Odrv4 I__256 (
            .O(N__1731),
            .I(\uart_tx.N_81 ));
    InMux I__255 (
            .O(N__1728),
            .I(N__1725));
    LocalMux I__254 (
            .O(N__1725),
            .I(\uart_tx.M_ctr_q_RNO_0Z0Z_2 ));
    InMux I__253 (
            .O(N__1722),
            .I(N__1718));
    InMux I__252 (
            .O(N__1721),
            .I(N__1715));
    LocalMux I__251 (
            .O(N__1718),
            .I(\uart_tx.M_ctr_qZ0Z_2 ));
    LocalMux I__250 (
            .O(N__1715),
            .I(\uart_tx.M_ctr_qZ0Z_2 ));
    CascadeMux I__249 (
            .O(N__1710),
            .I(\uart_rx.M_bitCtr_q_RNI578A4Z0Z_0_cascade_ ));
    InMux I__248 (
            .O(N__1707),
            .I(N__1702));
    InMux I__247 (
            .O(N__1706),
            .I(N__1699));
    InMux I__246 (
            .O(N__1705),
            .I(N__1696));
    LocalMux I__245 (
            .O(N__1702),
            .I(\uart_rx.M_ctr_qZ0Z_3 ));
    LocalMux I__244 (
            .O(N__1699),
            .I(\uart_rx.M_ctr_qZ0Z_3 ));
    LocalMux I__243 (
            .O(N__1696),
            .I(\uart_rx.M_ctr_qZ0Z_3 ));
    InMux I__242 (
            .O(N__1689),
            .I(N__1682));
    InMux I__241 (
            .O(N__1688),
            .I(N__1682));
    InMux I__240 (
            .O(N__1687),
            .I(N__1679));
    LocalMux I__239 (
            .O(N__1682),
            .I(\uart_rx.M_ctr_qZ0Z_5 ));
    LocalMux I__238 (
            .O(N__1679),
            .I(\uart_rx.M_ctr_qZ0Z_5 ));
    CascadeMux I__237 (
            .O(N__1674),
            .I(N__1671));
    InMux I__236 (
            .O(N__1671),
            .I(N__1665));
    InMux I__235 (
            .O(N__1670),
            .I(N__1660));
    InMux I__234 (
            .O(N__1669),
            .I(N__1660));
    InMux I__233 (
            .O(N__1668),
            .I(N__1657));
    LocalMux I__232 (
            .O(N__1665),
            .I(N__1654));
    LocalMux I__231 (
            .O(N__1660),
            .I(\uart_rx.M_ctr_qZ0Z_2 ));
    LocalMux I__230 (
            .O(N__1657),
            .I(\uart_rx.M_ctr_qZ0Z_2 ));
    Odrv4 I__229 (
            .O(N__1654),
            .I(\uart_rx.M_ctr_qZ0Z_2 ));
    InMux I__228 (
            .O(N__1647),
            .I(N__1642));
    InMux I__227 (
            .O(N__1646),
            .I(N__1637));
    InMux I__226 (
            .O(N__1645),
            .I(N__1637));
    LocalMux I__225 (
            .O(N__1642),
            .I(\uart_rx.M_ctr_qZ0Z_1 ));
    LocalMux I__224 (
            .O(N__1637),
            .I(\uart_rx.M_ctr_qZ0Z_1 ));
    InMux I__223 (
            .O(N__1632),
            .I(N__1629));
    LocalMux I__222 (
            .O(N__1629),
            .I(\uart_rx.M_ctr_q_RNIBJBV1Z0Z_1 ));
    CascadeMux I__221 (
            .O(N__1626),
            .I(N__1623));
    InMux I__220 (
            .O(N__1623),
            .I(N__1619));
    CascadeMux I__219 (
            .O(N__1622),
            .I(N__1616));
    LocalMux I__218 (
            .O(N__1619),
            .I(N__1612));
    InMux I__217 (
            .O(N__1616),
            .I(N__1607));
    InMux I__216 (
            .O(N__1615),
            .I(N__1607));
    Odrv4 I__215 (
            .O(N__1612),
            .I(\uart_rx.M_ctr_qZ0Z_6 ));
    LocalMux I__214 (
            .O(N__1607),
            .I(\uart_rx.M_ctr_qZ0Z_6 ));
    CascadeMux I__213 (
            .O(N__1602),
            .I(N__1599));
    InMux I__212 (
            .O(N__1599),
            .I(N__1593));
    InMux I__211 (
            .O(N__1598),
            .I(N__1590));
    InMux I__210 (
            .O(N__1597),
            .I(N__1587));
    InMux I__209 (
            .O(N__1596),
            .I(N__1584));
    LocalMux I__208 (
            .O(N__1593),
            .I(\uart_rx.M_ctr_qZ0Z_4 ));
    LocalMux I__207 (
            .O(N__1590),
            .I(\uart_rx.M_ctr_qZ0Z_4 ));
    LocalMux I__206 (
            .O(N__1587),
            .I(\uart_rx.M_ctr_qZ0Z_4 ));
    LocalMux I__205 (
            .O(N__1584),
            .I(\uart_rx.M_ctr_qZ0Z_4 ));
    CascadeMux I__204 (
            .O(N__1575),
            .I(\uart_rx.M_ctr_q_RNIBJBV1Z0Z_1_cascade_ ));
    InMux I__203 (
            .O(N__1572),
            .I(N__1563));
    InMux I__202 (
            .O(N__1571),
            .I(N__1563));
    InMux I__201 (
            .O(N__1570),
            .I(N__1556));
    InMux I__200 (
            .O(N__1569),
            .I(N__1556));
    InMux I__199 (
            .O(N__1568),
            .I(N__1556));
    LocalMux I__198 (
            .O(N__1563),
            .I(\uart_rx.M_ctr_qZ0Z_0 ));
    LocalMux I__197 (
            .O(N__1556),
            .I(\uart_rx.M_ctr_qZ0Z_0 ));
    CascadeMux I__196 (
            .O(N__1551),
            .I(\uart_rx.M_ctr_q_RNILBSE3Z0Z_6_cascade_ ));
    SRMux I__195 (
            .O(N__1548),
            .I(N__1545));
    LocalMux I__194 (
            .O(N__1545),
            .I(N__1542));
    Span4Mux_h I__193 (
            .O(N__1542),
            .I(N__1539));
    Span4Mux_s1_v I__192 (
            .O(N__1539),
            .I(N__1536));
    Odrv4 I__191 (
            .O(N__1536),
            .I(\uart_rx.M_state_q_RNIRDQO7_0Z0Z_0 ));
    CascadeMux I__190 (
            .O(N__1533),
            .I(uart_tx_N_187_1_cascade_));
    InMux I__189 (
            .O(N__1530),
            .I(N__1526));
    InMux I__188 (
            .O(N__1529),
            .I(N__1523));
    LocalMux I__187 (
            .O(N__1526),
            .I(\uart_tx.N_58 ));
    LocalMux I__186 (
            .O(N__1523),
            .I(\uart_tx.N_58 ));
    InMux I__185 (
            .O(N__1518),
            .I(N__1514));
    InMux I__184 (
            .O(N__1517),
            .I(N__1511));
    LocalMux I__183 (
            .O(N__1514),
            .I(\uart_tx.M_ctr_qZ0Z_3 ));
    LocalMux I__182 (
            .O(N__1511),
            .I(\uart_tx.M_ctr_qZ0Z_3 ));
    InMux I__181 (
            .O(N__1506),
            .I(\uart_tx.un1_M_ctr_q_3_cry_2 ));
    InMux I__180 (
            .O(N__1503),
            .I(N__1499));
    InMux I__179 (
            .O(N__1502),
            .I(N__1496));
    LocalMux I__178 (
            .O(N__1499),
            .I(\uart_tx.M_ctr_qZ0Z_4 ));
    LocalMux I__177 (
            .O(N__1496),
            .I(\uart_tx.M_ctr_qZ0Z_4 ));
    InMux I__176 (
            .O(N__1491),
            .I(\uart_tx.un1_M_ctr_q_3_cry_3 ));
    InMux I__175 (
            .O(N__1488),
            .I(\uart_tx.un1_M_ctr_q_3_cry_4 ));
    InMux I__174 (
            .O(N__1485),
            .I(\uart_tx.un1_M_ctr_q_3_cry_5 ));
    CascadeMux I__173 (
            .O(N__1482),
            .I(\uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_ ));
    CascadeMux I__172 (
            .O(N__1479),
            .I(N__1475));
    InMux I__171 (
            .O(N__1478),
            .I(N__1472));
    InMux I__170 (
            .O(N__1475),
            .I(N__1469));
    LocalMux I__169 (
            .O(N__1472),
            .I(\uart_tx.M_ctr_qZ0Z_6 ));
    LocalMux I__168 (
            .O(N__1469),
            .I(\uart_tx.M_ctr_qZ0Z_6 ));
    IoInMux I__167 (
            .O(N__1464),
            .I(N__1461));
    LocalMux I__166 (
            .O(N__1461),
            .I(usb_tx_c));
    InMux I__165 (
            .O(N__1458),
            .I(N__1455));
    LocalMux I__164 (
            .O(N__1455),
            .I(\uart_tx.M_txReg_d_0_iv_0_1 ));
    CascadeMux I__163 (
            .O(N__1452),
            .I(N__1449));
    InMux I__162 (
            .O(N__1449),
            .I(N__1439));
    InMux I__161 (
            .O(N__1448),
            .I(N__1439));
    InMux I__160 (
            .O(N__1447),
            .I(N__1439));
    InMux I__159 (
            .O(N__1446),
            .I(N__1436));
    LocalMux I__158 (
            .O(N__1439),
            .I(\uart_rx.un1_M_ctr_q_5_ac0_1_out ));
    LocalMux I__157 (
            .O(N__1436),
            .I(\uart_rx.un1_M_ctr_q_5_ac0_1_out ));
    CascadeMux I__156 (
            .O(N__1431),
            .I(\uart_tx.M_state_q_ns_0_o2_4_0_cascade_ ));
    CascadeMux I__155 (
            .O(N__1428),
            .I(\uart_tx.N_183_0_cascade_ ));
    CascadeMux I__154 (
            .O(N__1425),
            .I(\uart_tx.M_state_q_ns_0_i_0_0_0_cascade_ ));
    CascadeMux I__153 (
            .O(N__1422),
            .I(N__1418));
    InMux I__152 (
            .O(N__1421),
            .I(N__1415));
    InMux I__151 (
            .O(N__1418),
            .I(N__1412));
    LocalMux I__150 (
            .O(N__1415),
            .I(\uart_tx.N_187_1_i ));
    LocalMux I__149 (
            .O(N__1412),
            .I(\uart_tx.N_187_1_i ));
    InMux I__148 (
            .O(N__1407),
            .I(N__1403));
    InMux I__147 (
            .O(N__1406),
            .I(N__1400));
    LocalMux I__146 (
            .O(N__1403),
            .I(\uart_tx.M_ctr_qZ0Z_0 ));
    LocalMux I__145 (
            .O(N__1400),
            .I(\uart_tx.M_ctr_qZ0Z_0 ));
    InMux I__144 (
            .O(N__1395),
            .I(N__1391));
    InMux I__143 (
            .O(N__1394),
            .I(N__1388));
    LocalMux I__142 (
            .O(N__1391),
            .I(\uart_tx.M_ctr_qZ0Z_1 ));
    LocalMux I__141 (
            .O(N__1388),
            .I(\uart_tx.M_ctr_qZ0Z_1 ));
    InMux I__140 (
            .O(N__1383),
            .I(\uart_tx.un1_M_ctr_q_3_cry_0 ));
    InMux I__139 (
            .O(N__1380),
            .I(\uart_tx.un1_M_ctr_q_3_cry_1 ));
    CascadeMux I__138 (
            .O(N__1377),
            .I(\uart_rx.N_102_0_cascade_ ));
    CascadeMux I__137 (
            .O(N__1374),
            .I(N__1370));
    InMux I__136 (
            .O(N__1373),
            .I(N__1365));
    InMux I__135 (
            .O(N__1370),
            .I(N__1365));
    LocalMux I__134 (
            .O(N__1365),
            .I(\uart_rx.un1_M_ctr_q_5_ac0_7_0 ));
    InMux I__133 (
            .O(N__1362),
            .I(N__1344));
    InMux I__132 (
            .O(N__1361),
            .I(N__1344));
    InMux I__131 (
            .O(N__1360),
            .I(N__1344));
    InMux I__130 (
            .O(N__1359),
            .I(N__1344));
    InMux I__129 (
            .O(N__1358),
            .I(N__1344));
    InMux I__128 (
            .O(N__1357),
            .I(N__1344));
    LocalMux I__127 (
            .O(N__1344),
            .I(\uart_rx.N_102_0 ));
    InMux I__126 (
            .O(N__1341),
            .I(N__1338));
    LocalMux I__125 (
            .O(N__1338),
            .I(\uart_rx.un1_M_ctr_q_5_ac0_5_s_0_0 ));
    InMux I__124 (
            .O(N__1335),
            .I(N__1332));
    LocalMux I__123 (
            .O(N__1332),
            .I(\reset_cond.M_stage_qZ0Z_1 ));
    InMux I__122 (
            .O(N__1329),
            .I(N__1326));
    LocalMux I__121 (
            .O(N__1326),
            .I(\reset_cond.M_stage_qZ0Z_2 ));
    InMux I__120 (
            .O(N__1323),
            .I(N__1311));
    InMux I__119 (
            .O(N__1322),
            .I(N__1311));
    InMux I__118 (
            .O(N__1321),
            .I(N__1311));
    InMux I__117 (
            .O(N__1320),
            .I(N__1311));
    LocalMux I__116 (
            .O(N__1311),
            .I(N__1308));
    IoSpan4Mux I__115 (
            .O(N__1308),
            .I(N__1305));
    Odrv4 I__114 (
            .O(N__1305),
            .I(rst_n_c));
    InMux I__113 (
            .O(N__1302),
            .I(N__1299));
    LocalMux I__112 (
            .O(N__1299),
            .I(\reset_cond.M_stage_qZ0Z_0 ));
    CascadeMux I__111 (
            .O(N__1296),
            .I(\uart_rx.un1_M_ctr_q_5_ac0_5_s_0_0_cascade_ ));
    defparam IN_MUX_bfv_21_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_4_0_));
    defparam IN_MUX_bfv_23_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_23_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_23_4_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \reset_cond.M_stage_q_1_LC_20_2_0 .C_ON=1'b0;
    defparam \reset_cond.M_stage_q_1_LC_20_2_0 .SEQ_MODE=4'b1000;
    defparam \reset_cond.M_stage_q_1_LC_20_2_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \reset_cond.M_stage_q_1_LC_20_2_0  (
            .in0(N__1321),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1302),
            .lcout(\reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2539),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_cond.M_stage_q_2_LC_20_2_3 .C_ON=1'b0;
    defparam \reset_cond.M_stage_q_2_LC_20_2_3 .SEQ_MODE=4'b1000;
    defparam \reset_cond.M_stage_q_2_LC_20_2_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \reset_cond.M_stage_q_2_LC_20_2_3  (
            .in0(_gnd_net_),
            .in1(N__1322),
            .in2(_gnd_net_),
            .in3(N__1335),
            .lcout(\reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2539),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_cond.M_stage_q_3_LC_20_2_5 .C_ON=1'b0;
    defparam \reset_cond.M_stage_q_3_LC_20_2_5 .SEQ_MODE=4'b1000;
    defparam \reset_cond.M_stage_q_3_LC_20_2_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \reset_cond.M_stage_q_3_LC_20_2_5  (
            .in0(_gnd_net_),
            .in1(N__1323),
            .in2(_gnd_net_),
            .in3(N__1329),
            .lcout(M_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2539),
            .ce(),
            .sr(_gnd_net_));
    defparam \reset_cond.M_stage_q_0_LC_20_2_7 .C_ON=1'b0;
    defparam \reset_cond.M_stage_q_0_LC_20_2_7 .SEQ_MODE=4'b1000;
    defparam \reset_cond.M_stage_q_0_LC_20_2_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \reset_cond.M_stage_q_0_LC_20_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1320),
            .lcout(\reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2539),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_ctr_q_RNI5PLV_3_LC_21_1_4 .C_ON=1'b0;
    defparam \uart_rx.M_ctr_q_RNI5PLV_3_LC_21_1_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_ctr_q_RNI5PLV_3_LC_21_1_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_rx.M_ctr_q_RNI5PLV_3_LC_21_1_4  (
            .in0(_gnd_net_),
            .in1(N__1706),
            .in2(_gnd_net_),
            .in3(N__1668),
            .lcout(\uart_rx.un1_M_ctr_q_5_ac0_5_s_0_0 ),
            .ltout(\uart_rx.un1_M_ctr_q_5_ac0_5_s_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_ctr_q_RNIAC6F2_4_LC_21_1_5 .C_ON=1'b0;
    defparam \uart_rx.M_ctr_q_RNIAC6F2_4_LC_21_1_5 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_ctr_q_RNIAC6F2_4_LC_21_1_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \uart_rx.M_ctr_q_RNIAC6F2_4_LC_21_1_5  (
            .in0(_gnd_net_),
            .in1(N__1446),
            .in2(N__1296),
            .in3(N__1598),
            .lcout(\uart_rx.un1_M_ctr_q_5_ac0_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_ctr_q_0_LC_21_2_0 .C_ON=1'b0;
    defparam \uart_rx.M_ctr_q_0_LC_21_2_0 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_ctr_q_0_LC_21_2_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_rx.M_ctr_q_0_LC_21_2_0  (
            .in0(_gnd_net_),
            .in1(N__1571),
            .in2(_gnd_net_),
            .in3(N__1357),
            .lcout(\uart_rx.M_ctr_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2540),
            .ce(),
            .sr(N__1548));
    defparam \uart_rx.M_state_q_RNIRDQO7_0_LC_21_2_1 .C_ON=1'b0;
    defparam \uart_rx.M_state_q_RNIRDQO7_0_LC_21_2_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_state_q_RNIRDQO7_0_LC_21_2_1 .LUT_INIT=16'b0101100000001000;
    LogicCell40 \uart_rx.M_state_q_RNIRDQO7_0_LC_21_2_1  (
            .in0(N__2100),
            .in1(N__2169),
            .in2(N__2232),
            .in3(N__2329),
            .lcout(\uart_rx.N_102_0 ),
            .ltout(\uart_rx.N_102_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_ctr_q_1_LC_21_2_2 .C_ON=1'b0;
    defparam \uart_rx.M_ctr_q_1_LC_21_2_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_ctr_q_1_LC_21_2_2 .LUT_INIT=16'b0011111111000000;
    LogicCell40 \uart_rx.M_ctr_q_1_LC_21_2_2  (
            .in0(_gnd_net_),
            .in1(N__1572),
            .in2(N__1377),
            .in3(N__1647),
            .lcout(\uart_rx.M_ctr_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2540),
            .ce(),
            .sr(N__1548));
    defparam \uart_rx.M_ctr_q_5_LC_21_2_3 .C_ON=1'b0;
    defparam \uart_rx.M_ctr_q_5_LC_21_2_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_ctr_q_5_LC_21_2_3 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uart_rx.M_ctr_q_5_LC_21_2_3  (
            .in0(N__1360),
            .in1(_gnd_net_),
            .in2(N__1374),
            .in3(N__1689),
            .lcout(\uart_rx.M_ctr_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2540),
            .ce(),
            .sr(N__1548));
    defparam \uart_rx.M_ctr_q_6_LC_21_2_4 .C_ON=1'b0;
    defparam \uart_rx.M_ctr_q_6_LC_21_2_4 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_ctr_q_6_LC_21_2_4 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uart_rx.M_ctr_q_6_LC_21_2_4  (
            .in0(N__1688),
            .in1(N__1373),
            .in2(N__1626),
            .in3(N__1362),
            .lcout(\uart_rx.M_ctr_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2540),
            .ce(),
            .sr(N__1548));
    defparam \uart_rx.M_ctr_q_2_LC_21_2_5 .C_ON=1'b0;
    defparam \uart_rx.M_ctr_q_2_LC_21_2_5 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_ctr_q_2_LC_21_2_5 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uart_rx.M_ctr_q_2_LC_21_2_5  (
            .in0(N__1358),
            .in1(N__1447),
            .in2(_gnd_net_),
            .in3(N__1670),
            .lcout(\uart_rx.M_ctr_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2540),
            .ce(),
            .sr(N__1548));
    defparam \uart_rx.M_ctr_q_3_LC_21_2_6 .C_ON=1'b0;
    defparam \uart_rx.M_ctr_q_3_LC_21_2_6 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_ctr_q_3_LC_21_2_6 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uart_rx.M_ctr_q_3_LC_21_2_6  (
            .in0(N__1669),
            .in1(N__1361),
            .in2(N__1452),
            .in3(N__1707),
            .lcout(\uart_rx.M_ctr_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2540),
            .ce(),
            .sr(N__1548));
    defparam \uart_rx.M_ctr_q_4_LC_21_2_7 .C_ON=1'b0;
    defparam \uart_rx.M_ctr_q_4_LC_21_2_7 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_ctr_q_4_LC_21_2_7 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uart_rx.M_ctr_q_4_LC_21_2_7  (
            .in0(N__1359),
            .in1(N__1448),
            .in2(N__1602),
            .in3(N__1341),
            .lcout(\uart_rx.M_ctr_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2540),
            .ce(),
            .sr(N__1548));
    defparam \uart_tx.M_state_q_RNILEFM_0_LC_21_3_0 .C_ON=1'b0;
    defparam \uart_tx.M_state_q_RNILEFM_0_LC_21_3_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_state_q_RNILEFM_0_LC_21_3_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uart_tx.M_state_q_RNILEFM_0_LC_21_3_0  (
            .in0(_gnd_net_),
            .in1(N__1890),
            .in2(_gnd_net_),
            .in3(N__1819),
            .lcout(\uart_tx.N_187_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_state_q_RNILEFM_0_0_LC_21_3_1 .C_ON=1'b0;
    defparam \uart_tx.M_state_q_RNILEFM_0_0_LC_21_3_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_state_q_RNILEFM_0_0_LC_21_3_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uart_tx.M_state_q_RNILEFM_0_0_LC_21_3_1  (
            .in0(N__1820),
            .in1(_gnd_net_),
            .in2(N__1903),
            .in3(_gnd_net_),
            .lcout(\uart_tx.N_52_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_state_q_1_LC_21_3_2 .C_ON=1'b0;
    defparam \uart_tx.M_state_q_1_LC_21_3_2 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_state_q_1_LC_21_3_2 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uart_tx.M_state_q_1_LC_21_3_2  (
            .in0(N__2035),
            .in1(N__1895),
            .in2(N__1833),
            .in3(N__2139),
            .lcout(\uart_tx.M_state_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2542),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_RNIOOUF1_6_LC_21_3_3 .C_ON=1'b0;
    defparam \uart_tx.M_ctr_q_RNIOOUF1_6_LC_21_3_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_ctr_q_RNIOOUF1_6_LC_21_3_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uart_tx.M_ctr_q_RNIOOUF1_6_LC_21_3_3  (
            .in0(N__1965),
            .in1(N__1502),
            .in2(N__1479),
            .in3(N__1394),
            .lcout(),
            .ltout(\uart_tx.M_state_q_ns_0_o2_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_RNI3KTJ2_0_LC_21_3_4 .C_ON=1'b0;
    defparam \uart_tx.M_ctr_q_RNI3KTJ2_0_LC_21_3_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_ctr_q_RNI3KTJ2_0_LC_21_3_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uart_tx.M_ctr_q_RNI3KTJ2_0_LC_21_3_4  (
            .in0(N__1517),
            .in1(N__1722),
            .in2(N__1431),
            .in3(N__1407),
            .lcout(\uart_tx.N_183_0 ),
            .ltout(\uart_tx.N_183_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_bitCtr_q_RNIR97K3_1_LC_21_3_5 .C_ON=1'b0;
    defparam \uart_tx.M_bitCtr_q_RNIR97K3_1_LC_21_3_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_bitCtr_q_RNIR97K3_1_LC_21_3_5 .LUT_INIT=16'b1100111111111111;
    LogicCell40 \uart_tx.M_bitCtr_q_RNIR97K3_1_LC_21_3_5  (
            .in0(_gnd_net_),
            .in1(N__1866),
            .in2(N__1428),
            .in3(N__1765),
            .lcout(\uart_tx.N_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_state_q_RNO_0_0_LC_21_3_6 .C_ON=1'b0;
    defparam \uart_tx.M_state_q_RNO_0_0_LC_21_3_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_state_q_RNO_0_0_LC_21_3_6 .LUT_INIT=16'b0100010001110100;
    LogicCell40 \uart_tx.M_state_q_RNO_0_0_LC_21_3_6  (
            .in0(N__2034),
            .in1(N__1894),
            .in2(N__2984),
            .in3(N__1821),
            .lcout(),
            .ltout(\uart_tx.M_state_q_ns_0_i_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_state_q_0_LC_21_3_7 .C_ON=1'b0;
    defparam \uart_tx.M_state_q_0_LC_21_3_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_state_q_0_LC_21_3_7 .LUT_INIT=16'b0101000001010100;
    LogicCell40 \uart_tx.M_state_q_0_LC_21_3_7  (
            .in0(N__2138),
            .in1(N__2268),
            .in2(N__1425),
            .in3(N__1530),
            .lcout(\uart_tx.M_state_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2542),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_0_LC_21_4_0 .C_ON=1'b1;
    defparam \uart_tx.M_ctr_q_0_LC_21_4_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_0_LC_21_4_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \uart_tx.M_ctr_q_0_LC_21_4_0  (
            .in0(N__2870),
            .in1(N__1406),
            .in2(N__1422),
            .in3(N__1421),
            .lcout(\uart_tx.M_ctr_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_21_4_0_),
            .carryout(\uart_tx.un1_M_ctr_q_3_cry_0 ),
            .clk(N__2544),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_1_LC_21_4_1 .C_ON=1'b1;
    defparam \uart_tx.M_ctr_q_1_LC_21_4_1 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_1_LC_21_4_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \uart_tx.M_ctr_q_1_LC_21_4_1  (
            .in0(N__2874),
            .in1(N__1395),
            .in2(_gnd_net_),
            .in3(N__1383),
            .lcout(\uart_tx.M_ctr_qZ0Z_1 ),
            .ltout(),
            .carryin(\uart_tx.un1_M_ctr_q_3_cry_0 ),
            .carryout(\uart_tx.un1_M_ctr_q_3_cry_1 ),
            .clk(N__2544),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_RNO_0_2_LC_21_4_2 .C_ON=1'b1;
    defparam \uart_tx.M_ctr_q_RNO_0_2_LC_21_4_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_ctr_q_RNO_0_2_LC_21_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx.M_ctr_q_RNO_0_2_LC_21_4_2  (
            .in0(_gnd_net_),
            .in1(N__1721),
            .in2(_gnd_net_),
            .in3(N__1380),
            .lcout(\uart_tx.M_ctr_q_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\uart_tx.un1_M_ctr_q_3_cry_1 ),
            .carryout(\uart_tx.un1_M_ctr_q_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_3_LC_21_4_3 .C_ON=1'b1;
    defparam \uart_tx.M_ctr_q_3_LC_21_4_3 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_3_LC_21_4_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \uart_tx.M_ctr_q_3_LC_21_4_3  (
            .in0(N__2873),
            .in1(N__1518),
            .in2(_gnd_net_),
            .in3(N__1506),
            .lcout(\uart_tx.M_ctr_qZ0Z_3 ),
            .ltout(),
            .carryin(\uart_tx.un1_M_ctr_q_3_cry_2 ),
            .carryout(\uart_tx.un1_M_ctr_q_3_cry_3 ),
            .clk(N__2544),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_4_LC_21_4_4 .C_ON=1'b1;
    defparam \uart_tx.M_ctr_q_4_LC_21_4_4 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_4_LC_21_4_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \uart_tx.M_ctr_q_4_LC_21_4_4  (
            .in0(N__2871),
            .in1(N__1503),
            .in2(_gnd_net_),
            .in3(N__1491),
            .lcout(\uart_tx.M_ctr_qZ0Z_4 ),
            .ltout(),
            .carryin(\uart_tx.un1_M_ctr_q_3_cry_3 ),
            .carryout(\uart_tx.un1_M_ctr_q_3_cry_4 ),
            .clk(N__2544),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_RNO_0_5_LC_21_4_5 .C_ON=1'b1;
    defparam \uart_tx.M_ctr_q_RNO_0_5_LC_21_4_5 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_ctr_q_RNO_0_5_LC_21_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_tx.M_ctr_q_RNO_0_5_LC_21_4_5  (
            .in0(_gnd_net_),
            .in1(N__1964),
            .in2(_gnd_net_),
            .in3(N__1488),
            .lcout(\uart_tx.M_ctr_q_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\uart_tx.un1_M_ctr_q_3_cry_4 ),
            .carryout(\uart_tx.un1_M_ctr_q_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_RNO_0_6_LC_21_4_6 .C_ON=1'b0;
    defparam \uart_tx.M_ctr_q_RNO_0_6_LC_21_4_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_ctr_q_RNO_0_6_LC_21_4_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_tx.M_ctr_q_RNO_0_6_LC_21_4_6  (
            .in0(_gnd_net_),
            .in1(N__1478),
            .in2(_gnd_net_),
            .in3(N__1485),
            .lcout(),
            .ltout(\uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_6_LC_21_4_7 .C_ON=1'b0;
    defparam \uart_tx.M_ctr_q_6_LC_21_4_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_6_LC_21_4_7 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \uart_tx.M_ctr_q_6_LC_21_4_7  (
            .in0(N__1998),
            .in1(N__2872),
            .in2(N__1482),
            .in3(N__2038),
            .lcout(\uart_tx.M_ctr_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2544),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_txReg_q_LC_22_1_2 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_LC_22_1_2 .SEQ_MODE=4'b1001;
    defparam \uart_tx.M_txReg_q_LC_22_1_2 .LUT_INIT=16'b1110111110101111;
    LogicCell40 \uart_tx.M_txReg_q_LC_22_1_2  (
            .in0(N__1737),
            .in1(N__1458),
            .in2(N__2007),
            .in3(N__1832),
            .lcout(usb_tx_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2541),
            .ce(),
            .sr(N__2892));
    defparam \uart_tx.M_txReg_q_RNO_1_LC_22_2_0 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_RNO_1_LC_22_2_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_txReg_q_RNO_1_LC_22_2_0 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \uart_tx.M_txReg_q_RNO_1_LC_22_2_0  (
            .in0(N__1857),
            .in1(N__1911),
            .in2(N__2241),
            .in3(N__1770),
            .lcout(\uart_tx.M_txReg_d_0_iv_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_ctr_q_RNI1LLV_1_LC_22_2_1 .C_ON=1'b0;
    defparam \uart_rx.M_ctr_q_RNI1LLV_1_LC_22_2_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_ctr_q_RNI1LLV_1_LC_22_2_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_rx.M_ctr_q_RNI1LLV_1_LC_22_2_1  (
            .in0(N__1569),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1646),
            .lcout(\uart_rx.un1_M_ctr_q_5_ac0_1_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_state_q_ns_1_0__m19_0_o2_LC_22_2_2 .C_ON=1'b0;
    defparam \uart_rx.M_state_q_ns_1_0__m19_0_o2_LC_22_2_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_state_q_ns_1_0__m19_0_o2_LC_22_2_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \uart_rx.M_state_q_ns_1_0__m19_0_o2_LC_22_2_2  (
            .in0(N__1597),
            .in1(N__1570),
            .in2(N__1622),
            .in3(N__1632),
            .lcout(\uart_rx.m19_0_o2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_bitCtr_q_RNI578A4_0_LC_22_2_3 .C_ON=1'b0;
    defparam \uart_rx.M_bitCtr_q_RNI578A4_0_LC_22_2_3 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_bitCtr_q_RNI578A4_0_LC_22_2_3 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \uart_rx.M_bitCtr_q_RNI578A4_0_LC_22_2_3  (
            .in0(N__2090),
            .in1(N__2306),
            .in2(N__2226),
            .in3(N__2328),
            .lcout(\uart_rx.M_bitCtr_q_RNI578A4Z0Z_0 ),
            .ltout(\uart_rx.M_bitCtr_q_RNI578A4Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_state_q_ns_1_0__m19_0_a2_1_LC_22_2_4 .C_ON=1'b0;
    defparam \uart_rx.M_state_q_ns_1_0__m19_0_a2_1_LC_22_2_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_state_q_ns_1_0__m19_0_a2_1_LC_22_2_4 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \uart_rx.M_state_q_ns_1_0__m19_0_a2_1_LC_22_2_4  (
            .in0(N__2346),
            .in1(_gnd_net_),
            .in2(N__1710),
            .in3(N__1942),
            .lcout(\uart_rx.M_state_d_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_ctr_q_RNIBJBV1_1_LC_22_2_5 .C_ON=1'b0;
    defparam \uart_rx.M_ctr_q_RNIBJBV1_1_LC_22_2_5 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_ctr_q_RNIBJBV1_1_LC_22_2_5 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \uart_rx.M_ctr_q_RNIBJBV1_1_LC_22_2_5  (
            .in0(N__1705),
            .in1(N__1687),
            .in2(N__1674),
            .in3(N__1645),
            .lcout(\uart_rx.M_ctr_q_RNIBJBV1Z0Z_1 ),
            .ltout(\uart_rx.M_ctr_q_RNIBJBV1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_ctr_q_RNILBSE3_6_LC_22_2_6 .C_ON=1'b0;
    defparam \uart_rx.M_ctr_q_RNILBSE3_6_LC_22_2_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_ctr_q_RNILBSE3_6_LC_22_2_6 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \uart_rx.M_ctr_q_RNILBSE3_6_LC_22_2_6  (
            .in0(N__1615),
            .in1(N__1596),
            .in2(N__1575),
            .in3(N__1568),
            .lcout(\uart_rx.M_ctr_q_RNILBSE3Z0Z_6 ),
            .ltout(\uart_rx.M_ctr_q_RNILBSE3Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_state_q_RNIRDQO7_0_0_LC_22_2_7 .C_ON=1'b0;
    defparam \uart_rx.M_state_q_RNIRDQO7_0_0_LC_22_2_7 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_state_q_RNIRDQO7_0_0_LC_22_2_7 .LUT_INIT=16'b0001001101010111;
    LogicCell40 \uart_rx.M_state_q_RNIRDQO7_0_0_LC_22_2_7  (
            .in0(N__2212),
            .in1(N__2095),
            .in2(N__1551),
            .in3(N__2172),
            .lcout(\uart_rx.M_state_q_RNIRDQO7_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_0_LC_22_3_0 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_0_LC_22_3_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_0_LC_22_3_0 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \uart_tx.M_savedData_q_0_LC_22_3_0  (
            .in0(N__2046),
            .in1(N__2876),
            .in2(N__2977),
            .in3(N__1923),
            .lcout(\uart_tx.M_savedData_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2545),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_state_q_RNILEFM_1_0_LC_22_3_1 .C_ON=1'b0;
    defparam \uart_tx.M_state_q_RNILEFM_1_0_LC_22_3_1 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_state_q_RNILEFM_1_0_LC_22_3_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart_tx.M_state_q_RNILEFM_1_0_LC_22_3_1  (
            .in0(_gnd_net_),
            .in1(N__1896),
            .in2(_gnd_net_),
            .in3(N__1822),
            .lcout(uart_tx_N_187_1),
            .ltout(uart_tx_N_187_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_bitCtr_q_2_LC_22_3_2 .C_ON=1'b0;
    defparam \uart_tx.M_bitCtr_q_2_LC_22_3_2 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_bitCtr_q_2_LC_22_3_2 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \uart_tx.M_bitCtr_q_2_LC_22_3_2  (
            .in0(N__2265),
            .in1(_gnd_net_),
            .in2(N__1533),
            .in3(N__1529),
            .lcout(\uart_tx.M_bitCtr_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2545),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_txReg_q_RNO_5_LC_22_3_3 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_RNO_5_LC_22_3_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_txReg_q_RNO_5_LC_22_3_3 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \uart_tx.M_txReg_q_RNO_5_LC_22_3_3  (
            .in0(N__1922),
            .in1(N__2264),
            .in2(N__2499),
            .in3(N__1762),
            .lcout(),
            .ltout(\uart_tx.M_txReg_d_3_3_i_m4_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_txReg_q_RNO_4_LC_22_3_4 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_RNO_4_LC_22_3_4 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_txReg_q_RNO_4_LC_22_3_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \uart_tx.M_txReg_q_RNO_4_LC_22_3_4  (
            .in0(N__1763),
            .in1(N__2411),
            .in2(N__1914),
            .in3(N__2396),
            .lcout(\uart_tx.N_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_bitCtr_q_0_LC_22_3_5 .C_ON=1'b0;
    defparam \uart_tx.M_bitCtr_q_0_LC_22_3_5 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_bitCtr_q_0_LC_22_3_5 .LUT_INIT=16'b1111001000001000;
    LogicCell40 \uart_tx.M_bitCtr_q_0_LC_22_3_5  (
            .in0(N__1824),
            .in1(N__2037),
            .in2(N__1905),
            .in3(N__1852),
            .lcout(\uart_tx.M_bitCtr_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2545),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_bitCtr_q_RNIMHCR_0_LC_22_3_6 .C_ON=1'b0;
    defparam \uart_tx.M_bitCtr_q_RNIMHCR_0_LC_22_3_6 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_bitCtr_q_RNIMHCR_0_LC_22_3_6 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \uart_tx.M_bitCtr_q_RNIMHCR_0_LC_22_3_6  (
            .in0(N__1851),
            .in1(_gnd_net_),
            .in2(N__1904),
            .in3(N__1823),
            .lcout(\uart_tx.SUM_i_i_o4_1_1 ),
            .ltout(\uart_tx.SUM_i_i_o4_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_bitCtr_q_1_LC_22_3_7 .C_ON=1'b0;
    defparam \uart_tx.M_bitCtr_q_1_LC_22_3_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_bitCtr_q_1_LC_22_3_7 .LUT_INIT=16'b0101000100000100;
    LogicCell40 \uart_tx.M_bitCtr_q_1_LC_22_3_7  (
            .in0(N__2875),
            .in1(N__2036),
            .in2(N__1860),
            .in3(N__1764),
            .lcout(\uart_tx.M_bitCtr_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2545),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_3_LC_22_4_0 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_3_LC_22_4_0 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_3_LC_22_4_0 .LUT_INIT=16'b0010101011101010;
    LogicCell40 \uart_tx.M_savedData_q_3_LC_22_4_0  (
            .in0(N__1782),
            .in1(N__2879),
            .in2(N__2985),
            .in3(N__2373),
            .lcout(\uart_tx.M_savedData_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2548),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_txReg_q_RNO_2_LC_22_4_2 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_RNO_2_LC_22_4_2 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_txReg_q_RNO_2_LC_22_4_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_tx.M_txReg_q_RNO_2_LC_22_4_2  (
            .in0(_gnd_net_),
            .in1(N__1853),
            .in2(_gnd_net_),
            .in3(N__1825),
            .lcout(),
            .ltout(\uart_tx.M_txReg_d_0_iv_0_a2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_txReg_q_RNO_0_LC_22_4_3 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_RNO_0_LC_22_4_3 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_txReg_q_RNO_0_LC_22_4_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uart_tx.M_txReg_q_RNO_0_LC_22_4_3  (
            .in0(N__2267),
            .in1(N__1781),
            .in2(N__1773),
            .in3(N__1766),
            .lcout(\uart_tx.N_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_2_LC_22_4_5 .C_ON=1'b0;
    defparam \uart_tx.M_ctr_q_2_LC_22_4_5 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_2_LC_22_4_5 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \uart_tx.M_ctr_q_2_LC_22_4_5  (
            .in0(N__2877),
            .in1(N__2039),
            .in2(N__2002),
            .in3(N__1728),
            .lcout(\uart_tx.M_ctr_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2548),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_ctr_q_5_LC_22_4_7 .C_ON=1'b0;
    defparam \uart_tx.M_ctr_q_5_LC_22_4_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_ctr_q_5_LC_22_4_7 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \uart_tx.M_ctr_q_5_LC_22_4_7  (
            .in0(N__2878),
            .in1(N__2040),
            .in2(N__2003),
            .in3(N__1971),
            .lcout(\uart_tx.M_ctr_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2548),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.M_state_q_RNO_3_LC_23_1_1 .C_ON=1'b0;
    defparam \greeter.M_state_q_RNO_3_LC_23_1_1 .SEQ_MODE=4'b0000;
    defparam \greeter.M_state_q_RNO_3_LC_23_1_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \greeter.M_state_q_RNO_3_LC_23_1_1  (
            .in0(N__2426),
            .in1(N__3044),
            .in2(N__2484),
            .in3(N__3032),
            .lcout(),
            .ltout(\greeter.M_state_d_0_sqmuxa_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.M_state_q_RNO_1_LC_23_1_2 .C_ON=1'b0;
    defparam \greeter.M_state_q_RNO_1_LC_23_1_2 .SEQ_MODE=4'b0000;
    defparam \greeter.M_state_q_RNO_1_LC_23_1_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \greeter.M_state_q_RNO_1_LC_23_1_2  (
            .in0(N__2457),
            .in1(_gnd_net_),
            .in2(N__1950),
            .in3(N__2939),
            .lcout(\greeter.M_state_d_0_sqmuxa_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_state_q_ns_1_0__m22_0_LC_23_1_4 .C_ON=1'b0;
    defparam \uart_rx.M_state_q_ns_1_0__m22_0_LC_23_1_4 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_state_q_ns_1_0__m22_0_LC_23_1_4 .LUT_INIT=16'b0010101001101110;
    LogicCell40 \uart_rx.M_state_q_ns_1_0__m22_0_LC_23_1_4  (
            .in0(N__2208),
            .in1(N__2094),
            .in2(N__2584),
            .in3(N__2170),
            .lcout(),
            .ltout(\uart_rx.M_state_q_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_state_q_1_LC_23_1_5 .C_ON=1'b0;
    defparam \uart_rx.M_state_q_1_LC_23_1_5 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_state_q_1_LC_23_1_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \uart_rx.M_state_q_1_LC_23_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1947),
            .in3(N__2148),
            .lcout(\uart_rx.M_state_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2543),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_state_q_RNI62U94_0_LC_23_1_6 .C_ON=1'b0;
    defparam \uart_rx.M_state_q_RNI62U94_0_LC_23_1_6 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_state_q_RNI62U94_0_LC_23_1_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_rx.M_state_q_RNI62U94_0_LC_23_1_6  (
            .in0(N__2207),
            .in1(N__2093),
            .in2(_gnd_net_),
            .in3(N__2330),
            .lcout(\uart_rx.N_25_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_bitCtr_q_2_LC_23_2_0 .C_ON=1'b0;
    defparam \uart_rx.M_bitCtr_q_2_LC_23_2_0 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_bitCtr_q_2_LC_23_2_0 .LUT_INIT=16'b0010001100010000;
    LogicCell40 \uart_rx.M_bitCtr_q_2_LC_23_2_0  (
            .in0(N__2363),
            .in1(N__1929),
            .in2(N__2352),
            .in3(N__1943),
            .lcout(\uart_rx.M_bitCtr_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2546),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_newData_q_LC_23_2_1 .C_ON=1'b0;
    defparam \uart_rx.M_newData_q_LC_23_2_1 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_newData_q_LC_23_2_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_rx.M_newData_q_LC_23_2_1  (
            .in0(N__1944),
            .in1(N__2351),
            .in2(_gnd_net_),
            .in3(N__2364),
            .lcout(M_uart_rx_new_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2546),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_state_q_RNIHM1R_0_LC_23_2_2 .C_ON=1'b0;
    defparam \uart_rx.M_state_q_RNIHM1R_0_LC_23_2_2 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_state_q_RNIHM1R_0_LC_23_2_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart_rx.M_state_q_RNIHM1R_0_LC_23_2_2  (
            .in0(_gnd_net_),
            .in1(N__2216),
            .in2(_gnd_net_),
            .in3(N__2091),
            .lcout(\uart_rx.M_state_q_37_d ),
            .ltout(\uart_rx.M_state_q_37_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_bitCtr_q_1_LC_23_2_3 .C_ON=1'b0;
    defparam \uart_rx.M_bitCtr_q_1_LC_23_2_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_bitCtr_q_1_LC_23_2_3 .LUT_INIT=16'b0000110000000011;
    LogicCell40 \uart_rx.M_bitCtr_q_1_LC_23_2_3  (
            .in0(_gnd_net_),
            .in1(N__2347),
            .in2(N__2367),
            .in3(N__2362),
            .lcout(\uart_rx.M_bitCtr_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2546),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_bitCtr_q_0_LC_23_2_4 .C_ON=1'b0;
    defparam \uart_rx.M_bitCtr_q_0_LC_23_2_4 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_bitCtr_q_0_LC_23_2_4 .LUT_INIT=16'b1100100010011000;
    LogicCell40 \uart_rx.M_bitCtr_q_0_LC_23_2_4  (
            .in0(N__2092),
            .in1(N__2307),
            .in2(N__2228),
            .in3(N__2331),
            .lcout(\uart_rx.M_bitCtr_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2546),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.M_state_q_RNO_2_LC_23_2_5 .C_ON=1'b0;
    defparam \greeter.M_state_q_RNO_2_LC_23_2_5 .SEQ_MODE=4'b0000;
    defparam \greeter.M_state_q_RNO_2_LC_23_2_5 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \greeter.M_state_q_RNO_2_LC_23_2_5  (
            .in0(N__2940),
            .in1(N__2604),
            .in2(_gnd_net_),
            .in3(N__2859),
            .lcout(),
            .ltout(\greeter.M_state_q_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.M_state_q_LC_23_2_6 .C_ON=1'b0;
    defparam \greeter.M_state_q_LC_23_2_6 .SEQ_MODE=4'b1000;
    defparam \greeter.M_state_q_LC_23_2_6 .LUT_INIT=16'b0101010001010000;
    LogicCell40 \greeter.M_state_q_LC_23_2_6  (
            .in0(N__2140),
            .in1(N__2274),
            .in2(N__2295),
            .in3(N__2292),
            .lcout(greeter_M_state_q),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2546),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.M_state_q_RNO_0_LC_23_2_7 .C_ON=1'b0;
    defparam \greeter.M_state_q_RNO_0_LC_23_2_7 .SEQ_MODE=4'b0000;
    defparam \greeter.M_state_q_RNO_0_LC_23_2_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \greeter.M_state_q_RNO_0_LC_23_2_7  (
            .in0(N__2468),
            .in1(N__2450),
            .in2(N__2283),
            .in3(N__2438),
            .lcout(\greeter.M_state_d_0_sqmuxa_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_txReg_q_RNO_3_LC_23_3_0 .C_ON=1'b0;
    defparam \uart_tx.M_txReg_q_RNO_3_LC_23_3_0 .SEQ_MODE=4'b0000;
    defparam \uart_tx.M_txReg_q_RNO_3_LC_23_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart_tx.M_txReg_q_RNO_3_LC_23_3_0  (
            .in0(N__2996),
            .in1(N__2789),
            .in2(_gnd_net_),
            .in3(N__2266),
            .lcout(\uart_tx.N_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_state_q_ns_1_0__m19_0_0_LC_23_3_1 .C_ON=1'b0;
    defparam \uart_rx.M_state_q_ns_1_0__m19_0_0_LC_23_3_1 .SEQ_MODE=4'b0000;
    defparam \uart_rx.M_state_q_ns_1_0__m19_0_0_LC_23_3_1 .LUT_INIT=16'b0100110100001001;
    LogicCell40 \uart_rx.M_state_q_ns_1_0__m19_0_0_LC_23_3_1  (
            .in0(N__2227),
            .in1(N__2099),
            .in2(N__2589),
            .in3(N__2171),
            .lcout(),
            .ltout(\uart_rx.m19_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_state_q_0_LC_23_3_2 .C_ON=1'b0;
    defparam \uart_rx.M_state_q_0_LC_23_3_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_state_q_0_LC_23_3_2 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \uart_rx.M_state_q_0_LC_23_3_2  (
            .in0(N__2147),
            .in1(_gnd_net_),
            .in2(N__2109),
            .in3(N__2106),
            .lcout(\uart_rx.M_state_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2549),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.rom.letter_1_6_0__m5_0_LC_23_3_3 .C_ON=1'b0;
    defparam \greeter.rom.letter_1_6_0__m5_0_LC_23_3_3 .SEQ_MODE=4'b0000;
    defparam \greeter.rom.letter_1_6_0__m5_0_LC_23_3_3 .LUT_INIT=16'b0100101110000100;
    LogicCell40 \greeter.rom.letter_1_6_0__m5_0_LC_23_3_3  (
            .in0(N__2725),
            .in1(N__2638),
            .in2(N__2693),
            .in3(N__2764),
            .lcout(M_greeter_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.rom.letter_1_6_0__m23_i_LC_23_3_4 .C_ON=1'b0;
    defparam \greeter.rom.letter_1_6_0__m23_i_LC_23_3_4 .SEQ_MODE=4'b0000;
    defparam \greeter.rom.letter_1_6_0__m23_i_LC_23_3_4 .LUT_INIT=16'b1111100000100000;
    LogicCell40 \greeter.rom.letter_1_6_0__m23_i_LC_23_3_4  (
            .in0(N__2640),
            .in1(N__2727),
            .in2(N__2778),
            .in3(N__2684),
            .lcout(),
            .ltout(N_35_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_6_LC_23_3_5 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_6_LC_23_3_5 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_6_LC_23_3_5 .LUT_INIT=16'b0100111011001100;
    LogicCell40 \uart_tx.M_savedData_q_6_LC_23_3_5  (
            .in0(N__2960),
            .in1(N__2412),
            .in2(N__2415),
            .in3(N__2888),
            .lcout(\uart_tx.M_savedData_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2549),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.rom.letter_1_6_0__m12_i_LC_23_3_6 .C_ON=1'b0;
    defparam \greeter.rom.letter_1_6_0__m12_i_LC_23_3_6 .SEQ_MODE=4'b0000;
    defparam \greeter.rom.letter_1_6_0__m12_i_LC_23_3_6 .LUT_INIT=16'b1101100100100001;
    LogicCell40 \greeter.rom.letter_1_6_0__m12_i_LC_23_3_6  (
            .in0(N__2639),
            .in1(N__2726),
            .in2(N__2777),
            .in3(N__2683),
            .lcout(),
            .ltout(N_41_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_2_LC_23_3_7 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_2_LC_23_3_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_2_LC_23_3_7 .LUT_INIT=16'b0100111011001100;
    LogicCell40 \uart_tx.M_savedData_q_2_LC_23_3_7  (
            .in0(N__2959),
            .in1(N__2397),
            .in2(N__2400),
            .in3(N__2887),
            .lcout(\uart_tx.M_savedData_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2549),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.M_count_q_0_LC_23_4_0 .C_ON=1'b1;
    defparam \greeter.M_count_q_0_LC_23_4_0 .SEQ_MODE=4'b1000;
    defparam \greeter.M_count_q_0_LC_23_4_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \greeter.M_count_q_0_LC_23_4_0  (
            .in0(N__2972),
            .in1(N__2643),
            .in2(N__2884),
            .in3(N__2880),
            .lcout(\greeter.M_count_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_23_4_0_),
            .carryout(\greeter.un1_M_count_q_1_cry_0 ),
            .clk(N__2551),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.M_count_q_1_LC_23_4_1 .C_ON=1'b1;
    defparam \greeter.M_count_q_1_LC_23_4_1 .SEQ_MODE=4'b1000;
    defparam \greeter.M_count_q_1_LC_23_4_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \greeter.M_count_q_1_LC_23_4_1  (
            .in0(N__2975),
            .in1(N__2732),
            .in2(_gnd_net_),
            .in3(N__2382),
            .lcout(\greeter.M_count_qZ0Z_1 ),
            .ltout(),
            .carryin(\greeter.un1_M_count_q_1_cry_0 ),
            .carryout(\greeter.un1_M_count_q_1_cry_1 ),
            .clk(N__2551),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.M_count_q_2_LC_23_4_2 .C_ON=1'b1;
    defparam \greeter.M_count_q_2_LC_23_4_2 .SEQ_MODE=4'b1000;
    defparam \greeter.M_count_q_2_LC_23_4_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \greeter.M_count_q_2_LC_23_4_2  (
            .in0(N__2973),
            .in1(N__2773),
            .in2(_gnd_net_),
            .in3(N__2379),
            .lcout(\greeter.M_count_qZ1Z_2 ),
            .ltout(),
            .carryin(\greeter.un1_M_count_q_1_cry_1 ),
            .carryout(\greeter.un1_M_count_q_1_cry_2 ),
            .clk(N__2551),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.M_count_q_3_LC_23_4_3 .C_ON=1'b0;
    defparam \greeter.M_count_q_3_LC_23_4_3 .SEQ_MODE=4'b1000;
    defparam \greeter.M_count_q_3_LC_23_4_3 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \greeter.M_count_q_3_LC_23_4_3  (
            .in0(N__2689),
            .in1(N__2974),
            .in2(_gnd_net_),
            .in3(N__2376),
            .lcout(\greeter.M_count_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2551),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.rom.letter_1_6_0__m14_0_LC_23_4_5 .C_ON=1'b0;
    defparam \greeter.rom.letter_1_6_0__m14_0_LC_23_4_5 .SEQ_MODE=4'b0000;
    defparam \greeter.rom.letter_1_6_0__m14_0_LC_23_4_5 .LUT_INIT=16'b0100001101011000;
    LogicCell40 \greeter.rom.letter_1_6_0__m14_0_LC_23_4_5  (
            .in0(N__2771),
            .in1(N__2728),
            .in2(N__2694),
            .in3(N__2641),
            .lcout(m14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.rom.letter_1_6_0__m17_0_LC_23_4_6 .C_ON=1'b0;
    defparam \greeter.rom.letter_1_6_0__m17_0_LC_23_4_6 .SEQ_MODE=4'b0000;
    defparam \greeter.rom.letter_1_6_0__m17_0_LC_23_4_6 .LUT_INIT=16'b0001000000000100;
    LogicCell40 \greeter.rom.letter_1_6_0__m17_0_LC_23_4_6  (
            .in0(N__2642),
            .in1(N__2685),
            .in2(N__2733),
            .in3(N__2772),
            .lcout(),
            .ltout(M_greeter_tx_data_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_4_LC_23_4_7 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_4_LC_23_4_7 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_4_LC_23_4_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \uart_tx.M_savedData_q_4_LC_23_4_7  (
            .in0(N__2976),
            .in1(N__2858),
            .in2(N__2502),
            .in3(N__2498),
            .lcout(\uart_tx.M_savedData_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2551),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_savedData_q_6_LC_24_1_0 .C_ON=1'b0;
    defparam \uart_rx.M_savedData_q_6_LC_24_1_0 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_savedData_q_6_LC_24_1_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uart_rx.M_savedData_q_6_LC_24_1_0  (
            .in0(_gnd_net_),
            .in1(N__2483),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_uart_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2547),
            .ce(N__3017),
            .sr(_gnd_net_));
    defparam \uart_rx.M_savedData_q_7_LC_24_2_1 .C_ON=1'b0;
    defparam \uart_rx.M_savedData_q_7_LC_24_2_1 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_savedData_q_7_LC_24_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.M_savedData_q_7_LC_24_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2588),
            .lcout(M_uart_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2550),
            .ce(N__3021),
            .sr(_gnd_net_));
    defparam \uart_rx.M_savedData_q_2_LC_24_2_2 .C_ON=1'b0;
    defparam \uart_rx.M_savedData_q_2_LC_24_2_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_savedData_q_2_LC_24_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.M_savedData_q_2_LC_24_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3033),
            .lcout(M_uart_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2550),
            .ce(N__3021),
            .sr(_gnd_net_));
    defparam \uart_rx.M_savedData_q_5_LC_24_2_3 .C_ON=1'b0;
    defparam \uart_rx.M_savedData_q_5_LC_24_2_3 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_savedData_q_5_LC_24_2_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uart_rx.M_savedData_q_5_LC_24_2_3  (
            .in0(_gnd_net_),
            .in1(N__2469),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_uart_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2550),
            .ce(N__3021),
            .sr(_gnd_net_));
    defparam \uart_rx.M_savedData_q_0_LC_24_2_4 .C_ON=1'b0;
    defparam \uart_rx.M_savedData_q_0_LC_24_2_4 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_savedData_q_0_LC_24_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.M_savedData_q_0_LC_24_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2439),
            .lcout(M_uart_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2550),
            .ce(N__3021),
            .sr(_gnd_net_));
    defparam \uart_rx.M_savedData_q_1_LC_24_2_5 .C_ON=1'b0;
    defparam \uart_rx.M_savedData_q_1_LC_24_2_5 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_savedData_q_1_LC_24_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.M_savedData_q_1_LC_24_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2451),
            .lcout(M_uart_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2550),
            .ce(N__3021),
            .sr(_gnd_net_));
    defparam \uart_rx.M_savedData_q_4_LC_24_2_6 .C_ON=1'b0;
    defparam \uart_rx.M_savedData_q_4_LC_24_2_6 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_savedData_q_4_LC_24_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.M_savedData_q_4_LC_24_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2427),
            .lcout(M_uart_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2550),
            .ce(N__3021),
            .sr(_gnd_net_));
    defparam \uart_rx.M_savedData_q_3_LC_24_2_7 .C_ON=1'b0;
    defparam \uart_rx.M_savedData_q_3_LC_24_2_7 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_savedData_q_3_LC_24_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.M_savedData_q_3_LC_24_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3045),
            .lcout(M_uart_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2550),
            .ce(N__3021),
            .sr(_gnd_net_));
    defparam \greeter.rom.letter_1_6_0__m20_i_LC_24_3_2 .C_ON=1'b0;
    defparam \greeter.rom.letter_1_6_0__m20_i_LC_24_3_2 .SEQ_MODE=4'b0000;
    defparam \greeter.rom.letter_1_6_0__m20_i_LC_24_3_2 .LUT_INIT=16'b1010000010101001;
    LogicCell40 \greeter.rom.letter_1_6_0__m20_i_LC_24_3_2  (
            .in0(N__2775),
            .in1(N__2723),
            .in2(N__2691),
            .in3(N__2636),
            .lcout(),
            .ltout(N_37_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_5_LC_24_3_3 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_5_LC_24_3_3 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_5_LC_24_3_3 .LUT_INIT=16'b0100111011001100;
    LogicCell40 \uart_tx.M_savedData_q_5_LC_24_3_3  (
            .in0(N__2965),
            .in1(N__2997),
            .in2(N__3000),
            .in3(N__2886),
            .lcout(\uart_tx.M_savedData_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2552),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.rom.letter_1_6_0__m9_0_LC_24_3_4 .C_ON=1'b0;
    defparam \greeter.rom.letter_1_6_0__m9_0_LC_24_3_4 .SEQ_MODE=4'b0000;
    defparam \greeter.rom.letter_1_6_0__m9_0_LC_24_3_4 .LUT_INIT=16'b0000100000111010;
    LogicCell40 \greeter.rom.letter_1_6_0__m9_0_LC_24_3_4  (
            .in0(N__2776),
            .in1(N__2724),
            .in2(N__2692),
            .in3(N__2637),
            .lcout(),
            .ltout(M_greeter_tx_data_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_tx.M_savedData_q_1_LC_24_3_5 .C_ON=1'b0;
    defparam \uart_tx.M_savedData_q_1_LC_24_3_5 .SEQ_MODE=4'b1000;
    defparam \uart_tx.M_savedData_q_1_LC_24_3_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \uart_tx.M_savedData_q_1_LC_24_3_5  (
            .in0(N__2964),
            .in1(N__2790),
            .in2(N__2895),
            .in3(N__2885),
            .lcout(\uart_tx.M_savedData_qZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2552),
            .ce(),
            .sr(_gnd_net_));
    defparam \greeter.M_state_q_RNO_4_LC_24_3_6 .C_ON=1'b0;
    defparam \greeter.M_state_q_RNO_4_LC_24_3_6 .SEQ_MODE=4'b0000;
    defparam \greeter.M_state_q_RNO_4_LC_24_3_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \greeter.M_state_q_RNO_4_LC_24_3_6  (
            .in0(N__2774),
            .in1(N__2722),
            .in2(N__2690),
            .in3(N__2635),
            .lcout(\greeter.un1_M_state_d_0_sqmuxa_1_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_rx.M_rxd_q_LC_26_1_2 .C_ON=1'b0;
    defparam \uart_rx.M_rxd_q_LC_26_1_2 .SEQ_MODE=4'b1000;
    defparam \uart_rx.M_rxd_q_LC_26_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_rx.M_rxd_q_LC_26_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2598),
            .lcout(\uart_rx.M_rxd_qZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2553),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
