-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     Jun 12 2021 20:10:07

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    led : out std_logic_vector(7 downto 0);
    usb_tx : out std_logic;
    usb_rx : in std_logic;
    rst_n : in std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__3165\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2566\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2553\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2551\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2385\ : std_logic;
signal \N__2382\ : std_logic;
signal \N__2379\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2331\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2329\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2307\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2295\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2265\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2241\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2227\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2216\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2212\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2208\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2193\ : std_logic;
signal \N__2190\ : std_logic;
signal \N__2185\ : std_logic;
signal \N__2172\ : std_logic;
signal \N__2171\ : std_logic;
signal \N__2170\ : std_logic;
signal \N__2169\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2163\ : std_logic;
signal \N__2160\ : std_logic;
signal \N__2157\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2147\ : std_logic;
signal \N__2144\ : std_logic;
signal \N__2141\ : std_logic;
signal \N__2140\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2138\ : std_logic;
signal \N__2135\ : std_logic;
signal \N__2132\ : std_logic;
signal \N__2129\ : std_logic;
signal \N__2124\ : std_logic;
signal \N__2117\ : std_logic;
signal \N__2114\ : std_logic;
signal \N__2109\ : std_logic;
signal \N__2106\ : std_logic;
signal \N__2103\ : std_logic;
signal \N__2100\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2096\ : std_logic;
signal \N__2095\ : std_logic;
signal \N__2094\ : std_logic;
signal \N__2093\ : std_logic;
signal \N__2092\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2087\ : std_logic;
signal \N__2084\ : std_logic;
signal \N__2081\ : std_logic;
signal \N__2076\ : std_logic;
signal \N__2073\ : std_logic;
signal \N__2070\ : std_logic;
signal \N__2067\ : std_logic;
signal \N__2062\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2046\ : std_logic;
signal \N__2043\ : std_logic;
signal \N__2040\ : std_logic;
signal \N__2039\ : std_logic;
signal \N__2038\ : std_logic;
signal \N__2037\ : std_logic;
signal \N__2036\ : std_logic;
signal \N__2035\ : std_logic;
signal \N__2034\ : std_logic;
signal \N__2029\ : std_logic;
signal \N__2026\ : std_logic;
signal \N__2021\ : std_logic;
signal \N__2016\ : std_logic;
signal \N__2007\ : std_logic;
signal \N__2004\ : std_logic;
signal \N__2003\ : std_logic;
signal \N__2002\ : std_logic;
signal \N__1999\ : std_logic;
signal \N__1998\ : std_logic;
signal \N__1995\ : std_logic;
signal \N__1992\ : std_logic;
signal \N__1989\ : std_logic;
signal \N__1986\ : std_logic;
signal \N__1981\ : std_logic;
signal \N__1976\ : std_logic;
signal \N__1971\ : std_logic;
signal \N__1968\ : std_logic;
signal \N__1965\ : std_logic;
signal \N__1964\ : std_logic;
signal \N__1961\ : std_logic;
signal \N__1958\ : std_logic;
signal \N__1955\ : std_logic;
signal \N__1950\ : std_logic;
signal \N__1947\ : std_logic;
signal \N__1944\ : std_logic;
signal \N__1943\ : std_logic;
signal \N__1942\ : std_logic;
signal \N__1937\ : std_logic;
signal \N__1934\ : std_logic;
signal \N__1929\ : std_logic;
signal \N__1926\ : std_logic;
signal \N__1923\ : std_logic;
signal \N__1922\ : std_logic;
signal \N__1917\ : std_logic;
signal \N__1914\ : std_logic;
signal \N__1911\ : std_logic;
signal \N__1908\ : std_logic;
signal \N__1905\ : std_logic;
signal \N__1904\ : std_logic;
signal \N__1903\ : std_logic;
signal \N__1900\ : std_logic;
signal \N__1897\ : std_logic;
signal \N__1896\ : std_logic;
signal \N__1895\ : std_logic;
signal \N__1894\ : std_logic;
signal \N__1891\ : std_logic;
signal \N__1890\ : std_logic;
signal \N__1887\ : std_logic;
signal \N__1882\ : std_logic;
signal \N__1873\ : std_logic;
signal \N__1866\ : std_logic;
signal \N__1863\ : std_logic;
signal \N__1860\ : std_logic;
signal \N__1857\ : std_logic;
signal \N__1854\ : std_logic;
signal \N__1853\ : std_logic;
signal \N__1852\ : std_logic;
signal \N__1851\ : std_logic;
signal \N__1848\ : std_logic;
signal \N__1845\ : std_logic;
signal \N__1840\ : std_logic;
signal \N__1833\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1829\ : std_logic;
signal \N__1826\ : std_logic;
signal \N__1825\ : std_logic;
signal \N__1824\ : std_logic;
signal \N__1823\ : std_logic;
signal \N__1822\ : std_logic;
signal \N__1821\ : std_logic;
signal \N__1820\ : std_logic;
signal \N__1819\ : std_logic;
signal \N__1816\ : std_logic;
signal \N__1813\ : std_logic;
signal \N__1810\ : std_logic;
signal \N__1805\ : std_logic;
signal \N__1802\ : std_logic;
signal \N__1795\ : std_logic;
signal \N__1782\ : std_logic;
signal \N__1781\ : std_logic;
signal \N__1776\ : std_logic;
signal \N__1773\ : std_logic;
signal \N__1770\ : std_logic;
signal \N__1767\ : std_logic;
signal \N__1766\ : std_logic;
signal \N__1765\ : std_logic;
signal \N__1764\ : std_logic;
signal \N__1763\ : std_logic;
signal \N__1762\ : std_logic;
signal \N__1759\ : std_logic;
signal \N__1756\ : std_logic;
signal \N__1753\ : std_logic;
signal \N__1746\ : std_logic;
signal \N__1737\ : std_logic;
signal \N__1734\ : std_logic;
signal \N__1731\ : std_logic;
signal \N__1728\ : std_logic;
signal \N__1725\ : std_logic;
signal \N__1722\ : std_logic;
signal \N__1721\ : std_logic;
signal \N__1718\ : std_logic;
signal \N__1715\ : std_logic;
signal \N__1710\ : std_logic;
signal \N__1707\ : std_logic;
signal \N__1706\ : std_logic;
signal \N__1705\ : std_logic;
signal \N__1702\ : std_logic;
signal \N__1699\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1689\ : std_logic;
signal \N__1688\ : std_logic;
signal \N__1687\ : std_logic;
signal \N__1682\ : std_logic;
signal \N__1679\ : std_logic;
signal \N__1674\ : std_logic;
signal \N__1671\ : std_logic;
signal \N__1670\ : std_logic;
signal \N__1669\ : std_logic;
signal \N__1668\ : std_logic;
signal \N__1665\ : std_logic;
signal \N__1660\ : std_logic;
signal \N__1657\ : std_logic;
signal \N__1654\ : std_logic;
signal \N__1647\ : std_logic;
signal \N__1646\ : std_logic;
signal \N__1645\ : std_logic;
signal \N__1642\ : std_logic;
signal \N__1637\ : std_logic;
signal \N__1632\ : std_logic;
signal \N__1629\ : std_logic;
signal \N__1626\ : std_logic;
signal \N__1623\ : std_logic;
signal \N__1622\ : std_logic;
signal \N__1619\ : std_logic;
signal \N__1616\ : std_logic;
signal \N__1615\ : std_logic;
signal \N__1612\ : std_logic;
signal \N__1607\ : std_logic;
signal \N__1602\ : std_logic;
signal \N__1599\ : std_logic;
signal \N__1598\ : std_logic;
signal \N__1597\ : std_logic;
signal \N__1596\ : std_logic;
signal \N__1593\ : std_logic;
signal \N__1590\ : std_logic;
signal \N__1587\ : std_logic;
signal \N__1584\ : std_logic;
signal \N__1575\ : std_logic;
signal \N__1572\ : std_logic;
signal \N__1571\ : std_logic;
signal \N__1570\ : std_logic;
signal \N__1569\ : std_logic;
signal \N__1568\ : std_logic;
signal \N__1563\ : std_logic;
signal \N__1556\ : std_logic;
signal \N__1551\ : std_logic;
signal \N__1548\ : std_logic;
signal \N__1545\ : std_logic;
signal \N__1542\ : std_logic;
signal \N__1539\ : std_logic;
signal \N__1536\ : std_logic;
signal \N__1533\ : std_logic;
signal \N__1530\ : std_logic;
signal \N__1529\ : std_logic;
signal \N__1526\ : std_logic;
signal \N__1523\ : std_logic;
signal \N__1518\ : std_logic;
signal \N__1517\ : std_logic;
signal \N__1514\ : std_logic;
signal \N__1511\ : std_logic;
signal \N__1506\ : std_logic;
signal \N__1503\ : std_logic;
signal \N__1502\ : std_logic;
signal \N__1499\ : std_logic;
signal \N__1496\ : std_logic;
signal \N__1491\ : std_logic;
signal \N__1488\ : std_logic;
signal \N__1485\ : std_logic;
signal \N__1482\ : std_logic;
signal \N__1479\ : std_logic;
signal \N__1478\ : std_logic;
signal \N__1475\ : std_logic;
signal \N__1472\ : std_logic;
signal \N__1469\ : std_logic;
signal \N__1464\ : std_logic;
signal \N__1461\ : std_logic;
signal \N__1458\ : std_logic;
signal \N__1455\ : std_logic;
signal \N__1452\ : std_logic;
signal \N__1449\ : std_logic;
signal \N__1448\ : std_logic;
signal \N__1447\ : std_logic;
signal \N__1446\ : std_logic;
signal \N__1439\ : std_logic;
signal \N__1436\ : std_logic;
signal \N__1431\ : std_logic;
signal \N__1428\ : std_logic;
signal \N__1425\ : std_logic;
signal \N__1422\ : std_logic;
signal \N__1421\ : std_logic;
signal \N__1418\ : std_logic;
signal \N__1415\ : std_logic;
signal \N__1412\ : std_logic;
signal \N__1407\ : std_logic;
signal \N__1406\ : std_logic;
signal \N__1403\ : std_logic;
signal \N__1400\ : std_logic;
signal \N__1395\ : std_logic;
signal \N__1394\ : std_logic;
signal \N__1391\ : std_logic;
signal \N__1388\ : std_logic;
signal \N__1383\ : std_logic;
signal \N__1380\ : std_logic;
signal \N__1377\ : std_logic;
signal \N__1374\ : std_logic;
signal \N__1373\ : std_logic;
signal \N__1370\ : std_logic;
signal \N__1365\ : std_logic;
signal \N__1362\ : std_logic;
signal \N__1361\ : std_logic;
signal \N__1360\ : std_logic;
signal \N__1359\ : std_logic;
signal \N__1358\ : std_logic;
signal \N__1357\ : std_logic;
signal \N__1344\ : std_logic;
signal \N__1341\ : std_logic;
signal \N__1338\ : std_logic;
signal \N__1335\ : std_logic;
signal \N__1332\ : std_logic;
signal \N__1329\ : std_logic;
signal \N__1326\ : std_logic;
signal \N__1323\ : std_logic;
signal \N__1322\ : std_logic;
signal \N__1321\ : std_logic;
signal \N__1320\ : std_logic;
signal \N__1311\ : std_logic;
signal \N__1308\ : std_logic;
signal \N__1305\ : std_logic;
signal \N__1302\ : std_logic;
signal \N__1299\ : std_logic;
signal \N__1296\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal rst_n_c : std_logic;
signal \reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \uart_rx.un1_M_ctr_q_5_ac0_5_s_0_0_cascade_\ : std_logic;
signal \uart_rx.N_102_0_cascade_\ : std_logic;
signal \uart_rx.un1_M_ctr_q_5_ac0_7_0\ : std_logic;
signal \uart_rx.N_102_0\ : std_logic;
signal \uart_rx.un1_M_ctr_q_5_ac0_5_s_0_0\ : std_logic;
signal \uart_tx.M_state_q_ns_0_o2_4_0_cascade_\ : std_logic;
signal \uart_tx.N_183_0_cascade_\ : std_logic;
signal \uart_tx.M_state_q_ns_0_i_0_0_0_cascade_\ : std_logic;
signal \uart_tx.N_187_1_i\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_0\ : std_logic;
signal \bfn_21_4_0_\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_1\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_0\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_1\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_3\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_2\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_4\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_3\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_4\ : std_logic;
signal \uart_tx.un1_M_ctr_q_3_cry_5\ : std_logic;
signal \uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_6\ : std_logic;
signal usb_tx_c : std_logic;
signal \uart_tx.M_txReg_d_0_iv_0_1\ : std_logic;
signal \uart_rx.un1_M_ctr_q_5_ac0_1_out\ : std_logic;
signal \uart_rx.M_bitCtr_q_RNI578A4Z0Z_0_cascade_\ : std_logic;
signal \uart_rx.M_ctr_qZ0Z_3\ : std_logic;
signal \uart_rx.M_ctr_qZ0Z_5\ : std_logic;
signal \uart_rx.M_ctr_qZ0Z_2\ : std_logic;
signal \uart_rx.M_ctr_qZ0Z_1\ : std_logic;
signal \uart_rx.M_ctr_q_RNIBJBV1Z0Z_1\ : std_logic;
signal \uart_rx.M_ctr_qZ0Z_6\ : std_logic;
signal \uart_rx.M_ctr_qZ0Z_4\ : std_logic;
signal \uart_rx.M_ctr_q_RNIBJBV1Z0Z_1_cascade_\ : std_logic;
signal \uart_rx.M_ctr_qZ0Z_0\ : std_logic;
signal \uart_rx.M_ctr_q_RNILBSE3Z0Z_6_cascade_\ : std_logic;
signal \uart_rx.M_state_q_RNIRDQO7_0Z0Z_0\ : std_logic;
signal \uart_tx_N_187_1_cascade_\ : std_logic;
signal \uart_tx.N_58\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_0\ : std_logic;
signal \uart_tx.M_txReg_d_3_3_i_m4_ns_1_cascade_\ : std_logic;
signal \uart_tx.N_66\ : std_logic;
signal \uart_tx.M_state_qZ0Z_0\ : std_logic;
signal \uart_tx.SUM_i_i_o4_1_1\ : std_logic;
signal \uart_tx.SUM_i_i_o4_1_1_cascade_\ : std_logic;
signal \uart_tx.M_bitCtr_qZ0Z_0\ : std_logic;
signal \uart_tx.M_state_qZ0Z_1\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_3\ : std_logic;
signal \uart_tx.M_txReg_d_0_iv_0_a2_1_1_cascade_\ : std_logic;
signal \uart_tx.M_bitCtr_qZ0Z_1\ : std_logic;
signal \uart_tx.N_81\ : std_logic;
signal \uart_tx.M_ctr_q_RNO_0Z0Z_2\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_2\ : std_logic;
signal \uart_tx.N_183_0\ : std_logic;
signal \uart_tx.N_52_i\ : std_logic;
signal \uart_tx.M_ctr_q_RNO_0Z0Z_5\ : std_logic;
signal \uart_tx.M_ctr_qZ0Z_5\ : std_logic;
signal \greeter.M_state_d_0_sqmuxa_1_5_cascade_\ : std_logic;
signal \uart_rx.M_state_q_ns_1_cascade_\ : std_logic;
signal \uart_rx.M_bitCtr_qZ0Z_2\ : std_logic;
signal \uart_rx.M_state_q_37_d\ : std_logic;
signal \uart_rx.M_state_q_37_d_cascade_\ : std_logic;
signal \uart_rx.M_bitCtr_q_RNI578A4Z0Z_0\ : std_logic;
signal \uart_rx.M_bitCtr_qZ0Z_1\ : std_logic;
signal \uart_rx.M_ctr_q_RNILBSE3Z0Z_6\ : std_logic;
signal \uart_rx.M_bitCtr_qZ0Z_0\ : std_logic;
signal \greeter.M_state_q_0_cascade_\ : std_logic;
signal \greeter.M_state_d_0_sqmuxa_1_7\ : std_logic;
signal \M_uart_rx_new_data_0\ : std_logic;
signal \greeter.M_state_d_0_sqmuxa_1_6\ : std_logic;
signal \uart_tx.M_bitCtr_qZ0Z_2\ : std_logic;
signal \uart_tx.N_65\ : std_logic;
signal \uart_rx.M_state_qZ0Z_1\ : std_logic;
signal \uart_rx.m19_0_o2\ : std_logic;
signal \M_reset_cond_out_0\ : std_logic;
signal \uart_rx.m19_0_0_cascade_\ : std_logic;
signal \uart_rx.M_state_d_0_sqmuxa_1\ : std_logic;
signal \uart_rx.M_state_qZ0Z_0\ : std_logic;
signal \M_greeter_tx_data_0\ : std_logic;
signal \N_35_cascade_\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_6\ : std_logic;
signal \N_41_cascade_\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_2\ : std_logic;
signal \bfn_23_4_0_\ : std_logic;
signal \greeter.un1_M_count_q_1_cry_0\ : std_logic;
signal \greeter.un1_M_count_q_1_cry_1\ : std_logic;
signal \greeter.un1_M_count_q_1_cry_2\ : std_logic;
signal m14_0 : std_logic;
signal \M_greeter_tx_data_4_cascade_\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_4\ : std_logic;
signal \M_uart_rx_data_7\ : std_logic;
signal \M_uart_rx_data_6\ : std_logic;
signal \M_uart_rx_data_0\ : std_logic;
signal \M_uart_rx_data_2\ : std_logic;
signal \M_uart_rx_data_1\ : std_logic;
signal \M_uart_rx_data_5\ : std_logic;
signal \M_uart_rx_data_4\ : std_logic;
signal \M_uart_rx_data_3\ : std_logic;
signal \uart_rx.N_25_i\ : std_logic;
signal \N_37_cascade_\ : std_logic;
signal \uart_tx.M_savedData_qZ0Z_5\ : std_logic;
signal \greeter_M_state_q\ : std_logic;
signal \M_greeter_tx_data_1_cascade_\ : std_logic;
signal \uart_tx_N_187_1\ : std_logic;
signal \uart_tx.M_savedData_qZ1Z_1\ : std_logic;
signal \greeter.M_count_qZ1Z_2\ : std_logic;
signal \greeter.M_count_qZ0Z_1\ : std_logic;
signal \greeter.M_count_qZ0Z_3\ : std_logic;
signal \greeter.M_count_qZ0Z_0\ : std_logic;
signal \greeter.un1_M_state_d_0_sqmuxa_1_0_a2_0_0\ : std_logic;
signal usb_rx_c : std_logic;
signal \uart_rx.M_rxd_qZ0\ : std_logic;
signal clk_c_g : std_logic;
signal \_gnd_net_\ : std_logic;

signal clk_wire : std_logic;
signal led_wire : std_logic_vector(7 downto 0);
signal rst_n_wire : std_logic;
signal usb_rx_wire : std_logic;
signal usb_tx_wire : std_logic;

begin
    clk_wire <= clk;
    led <= led_wire;
    rst_n_wire <= rst_n;
    usb_rx_wire <= usb_rx;
    usb_tx <= usb_tx_wire;

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__3163\,
            GLOBALBUFFEROUTPUT => clk_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3165\,
            DIN => \N__3164\,
            DOUT => \N__3163\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3165\,
            PADOUT => \N__3164\,
            PADIN => \N__3163\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3154\,
            DIN => \N__3153\,
            DOUT => \N__3152\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3154\,
            PADOUT => \N__3153\,
            PADIN => \N__3152\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3145\,
            DIN => \N__3144\,
            DOUT => \N__3143\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3145\,
            PADOUT => \N__3144\,
            PADIN => \N__3143\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3136\,
            DIN => \N__3135\,
            DOUT => \N__3134\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3136\,
            PADOUT => \N__3135\,
            PADIN => \N__3134\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3127\,
            DIN => \N__3126\,
            DOUT => \N__3125\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3127\,
            PADOUT => \N__3126\,
            PADIN => \N__3125\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3118\,
            DIN => \N__3117\,
            DOUT => \N__3116\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3118\,
            PADOUT => \N__3117\,
            PADIN => \N__3116\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3109\,
            DIN => \N__3108\,
            DOUT => \N__3107\,
            PACKAGEPIN => led_wire(5)
        );

    \led_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3109\,
            PADOUT => \N__3108\,
            PADIN => \N__3107\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3100\,
            DIN => \N__3099\,
            DOUT => \N__3098\,
            PACKAGEPIN => led_wire(6)
        );

    \led_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3100\,
            PADOUT => \N__3099\,
            PADIN => \N__3098\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3091\,
            DIN => \N__3090\,
            DOUT => \N__3089\,
            PACKAGEPIN => led_wire(7)
        );

    \led_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3091\,
            PADOUT => \N__3090\,
            PADIN => \N__3089\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3082\,
            DIN => \N__3081\,
            DOUT => \N__3080\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3082\,
            PADOUT => \N__3081\,
            PADIN => \N__3080\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \usb_rx_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3073\,
            DIN => \N__3072\,
            DOUT => \N__3071\,
            PACKAGEPIN => usb_rx_wire
        );

    \usb_rx_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3073\,
            PADOUT => \N__3072\,
            PADIN => \N__3071\,
            CLOCKENABLE => 'H',
            DIN0 => usb_rx_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \usb_tx_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3064\,
            DIN => \N__3063\,
            DOUT => \N__3062\,
            PACKAGEPIN => usb_tx_wire
        );

    \usb_tx_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3064\,
            PADOUT => \N__3063\,
            PADIN => \N__3062\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1464\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__694\ : InMux
    port map (
            O => \N__3045\,
            I => \N__3041\
        );

    \I__693\ : InMux
    port map (
            O => \N__3044\,
            I => \N__3038\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__3041\,
            I => \M_uart_rx_data_4\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__3038\,
            I => \M_uart_rx_data_4\
        );

    \I__690\ : InMux
    port map (
            O => \N__3033\,
            I => \N__3029\
        );

    \I__689\ : InMux
    port map (
            O => \N__3032\,
            I => \N__3026\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3029\,
            I => \M_uart_rx_data_3\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3026\,
            I => \M_uart_rx_data_3\
        );

    \I__686\ : CEMux
    port map (
            O => \N__3021\,
            I => \N__3018\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__3018\,
            I => \N__3014\
        );

    \I__684\ : CEMux
    port map (
            O => \N__3017\,
            I => \N__3011\
        );

    \I__683\ : Span4Mux_v
    port map (
            O => \N__3014\,
            I => \N__3006\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__3011\,
            I => \N__3006\
        );

    \I__681\ : Span4Mux_s0_v
    port map (
            O => \N__3006\,
            I => \N__3003\
        );

    \I__680\ : Odrv4
    port map (
            O => \N__3003\,
            I => \uart_rx.N_25_i\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__3000\,
            I => \N_37_cascade_\
        );

    \I__678\ : InMux
    port map (
            O => \N__2997\,
            I => \N__2993\
        );

    \I__677\ : InMux
    port map (
            O => \N__2996\,
            I => \N__2990\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__2993\,
            I => \uart_tx.M_savedData_qZ0Z_5\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__2990\,
            I => \uart_tx.M_savedData_qZ0Z_5\
        );

    \I__674\ : CascadeMux
    port map (
            O => \N__2985\,
            I => \N__2981\
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__2984\,
            I => \N__2978\
        );

    \I__672\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2969\
        );

    \I__671\ : InMux
    port map (
            O => \N__2978\,
            I => \N__2966\
        );

    \I__670\ : CascadeMux
    port map (
            O => \N__2977\,
            I => \N__2961\
        );

    \I__669\ : InMux
    port map (
            O => \N__2976\,
            I => \N__2954\
        );

    \I__668\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2954\
        );

    \I__667\ : InMux
    port map (
            O => \N__2974\,
            I => \N__2947\
        );

    \I__666\ : InMux
    port map (
            O => \N__2973\,
            I => \N__2947\
        );

    \I__665\ : InMux
    port map (
            O => \N__2972\,
            I => \N__2947\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__2969\,
            I => \N__2944\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__2966\,
            I => \N__2941\
        );

    \I__662\ : InMux
    port map (
            O => \N__2965\,
            I => \N__2934\
        );

    \I__661\ : InMux
    port map (
            O => \N__2964\,
            I => \N__2934\
        );

    \I__660\ : InMux
    port map (
            O => \N__2961\,
            I => \N__2931\
        );

    \I__659\ : InMux
    port map (
            O => \N__2960\,
            I => \N__2926\
        );

    \I__658\ : InMux
    port map (
            O => \N__2959\,
            I => \N__2926\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__2954\,
            I => \N__2921\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__2947\,
            I => \N__2921\
        );

    \I__655\ : Span4Mux_v
    port map (
            O => \N__2944\,
            I => \N__2916\
        );

    \I__654\ : Span4Mux_h
    port map (
            O => \N__2941\,
            I => \N__2916\
        );

    \I__653\ : InMux
    port map (
            O => \N__2940\,
            I => \N__2913\
        );

    \I__652\ : InMux
    port map (
            O => \N__2939\,
            I => \N__2910\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__2934\,
            I => \greeter_M_state_q\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__2931\,
            I => \greeter_M_state_q\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__2926\,
            I => \greeter_M_state_q\
        );

    \I__648\ : Odrv4
    port map (
            O => \N__2921\,
            I => \greeter_M_state_q\
        );

    \I__647\ : Odrv4
    port map (
            O => \N__2916\,
            I => \greeter_M_state_q\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__2913\,
            I => \greeter_M_state_q\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__2910\,
            I => \greeter_M_state_q\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__2895\,
            I => \M_greeter_tx_data_1_cascade_\
        );

    \I__643\ : SRMux
    port map (
            O => \N__2892\,
            I => \N__2889\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__2889\,
            I => \N__2881\
        );

    \I__641\ : InMux
    port map (
            O => \N__2888\,
            I => \N__2865\
        );

    \I__640\ : InMux
    port map (
            O => \N__2887\,
            I => \N__2865\
        );

    \I__639\ : InMux
    port map (
            O => \N__2886\,
            I => \N__2860\
        );

    \I__638\ : InMux
    port map (
            O => \N__2885\,
            I => \N__2860\
        );

    \I__637\ : CascadeMux
    port map (
            O => \N__2884\,
            I => \N__2855\
        );

    \I__636\ : Span4Mux_h
    port map (
            O => \N__2881\,
            I => \N__2852\
        );

    \I__635\ : InMux
    port map (
            O => \N__2880\,
            I => \N__2849\
        );

    \I__634\ : InMux
    port map (
            O => \N__2879\,
            I => \N__2842\
        );

    \I__633\ : InMux
    port map (
            O => \N__2878\,
            I => \N__2842\
        );

    \I__632\ : InMux
    port map (
            O => \N__2877\,
            I => \N__2842\
        );

    \I__631\ : InMux
    port map (
            O => \N__2876\,
            I => \N__2837\
        );

    \I__630\ : InMux
    port map (
            O => \N__2875\,
            I => \N__2837\
        );

    \I__629\ : InMux
    port map (
            O => \N__2874\,
            I => \N__2832\
        );

    \I__628\ : InMux
    port map (
            O => \N__2873\,
            I => \N__2832\
        );

    \I__627\ : InMux
    port map (
            O => \N__2872\,
            I => \N__2825\
        );

    \I__626\ : InMux
    port map (
            O => \N__2871\,
            I => \N__2825\
        );

    \I__625\ : InMux
    port map (
            O => \N__2870\,
            I => \N__2825\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__2865\,
            I => \N__2820\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__2860\,
            I => \N__2820\
        );

    \I__622\ : InMux
    port map (
            O => \N__2859\,
            I => \N__2817\
        );

    \I__621\ : InMux
    port map (
            O => \N__2858\,
            I => \N__2812\
        );

    \I__620\ : InMux
    port map (
            O => \N__2855\,
            I => \N__2812\
        );

    \I__619\ : Span4Mux_s0_v
    port map (
            O => \N__2852\,
            I => \N__2809\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__2849\,
            I => \uart_tx_N_187_1\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__2842\,
            I => \uart_tx_N_187_1\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__2837\,
            I => \uart_tx_N_187_1\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__2832\,
            I => \uart_tx_N_187_1\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__2825\,
            I => \uart_tx_N_187_1\
        );

    \I__613\ : Odrv4
    port map (
            O => \N__2820\,
            I => \uart_tx_N_187_1\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__2817\,
            I => \uart_tx_N_187_1\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__2812\,
            I => \uart_tx_N_187_1\
        );

    \I__610\ : Odrv4
    port map (
            O => \N__2809\,
            I => \uart_tx_N_187_1\
        );

    \I__609\ : InMux
    port map (
            O => \N__2790\,
            I => \N__2786\
        );

    \I__608\ : InMux
    port map (
            O => \N__2789\,
            I => \N__2783\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__2786\,
            I => \uart_tx.M_savedData_qZ1Z_1\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__2783\,
            I => \uart_tx.M_savedData_qZ1Z_1\
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__2778\,
            I => \N__2768\
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__2777\,
            I => \N__2765\
        );

    \I__603\ : InMux
    port map (
            O => \N__2776\,
            I => \N__2757\
        );

    \I__602\ : InMux
    port map (
            O => \N__2775\,
            I => \N__2757\
        );

    \I__601\ : InMux
    port map (
            O => \N__2774\,
            I => \N__2757\
        );

    \I__600\ : InMux
    port map (
            O => \N__2773\,
            I => \N__2750\
        );

    \I__599\ : InMux
    port map (
            O => \N__2772\,
            I => \N__2750\
        );

    \I__598\ : InMux
    port map (
            O => \N__2771\,
            I => \N__2750\
        );

    \I__597\ : InMux
    port map (
            O => \N__2768\,
            I => \N__2743\
        );

    \I__596\ : InMux
    port map (
            O => \N__2765\,
            I => \N__2743\
        );

    \I__595\ : InMux
    port map (
            O => \N__2764\,
            I => \N__2743\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__2757\,
            I => \N__2740\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__2750\,
            I => \greeter.M_count_qZ1Z_2\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__2743\,
            I => \greeter.M_count_qZ1Z_2\
        );

    \I__591\ : Odrv4
    port map (
            O => \N__2740\,
            I => \greeter.M_count_qZ1Z_2\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__2733\,
            I => \N__2729\
        );

    \I__589\ : InMux
    port map (
            O => \N__2732\,
            I => \N__2715\
        );

    \I__588\ : InMux
    port map (
            O => \N__2729\,
            I => \N__2715\
        );

    \I__587\ : InMux
    port map (
            O => \N__2728\,
            I => \N__2715\
        );

    \I__586\ : InMux
    port map (
            O => \N__2727\,
            I => \N__2708\
        );

    \I__585\ : InMux
    port map (
            O => \N__2726\,
            I => \N__2708\
        );

    \I__584\ : InMux
    port map (
            O => \N__2725\,
            I => \N__2708\
        );

    \I__583\ : InMux
    port map (
            O => \N__2724\,
            I => \N__2701\
        );

    \I__582\ : InMux
    port map (
            O => \N__2723\,
            I => \N__2701\
        );

    \I__581\ : InMux
    port map (
            O => \N__2722\,
            I => \N__2701\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__2715\,
            I => \greeter.M_count_qZ0Z_1\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__2708\,
            I => \greeter.M_count_qZ0Z_1\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__2701\,
            I => \greeter.M_count_qZ0Z_1\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__2694\,
            I => \N__2686\
        );

    \I__576\ : CascadeMux
    port map (
            O => \N__2693\,
            I => \N__2680\
        );

    \I__575\ : CascadeMux
    port map (
            O => \N__2692\,
            I => \N__2677\
        );

    \I__574\ : CascadeMux
    port map (
            O => \N__2691\,
            I => \N__2674\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__2690\,
            I => \N__2671\
        );

    \I__572\ : InMux
    port map (
            O => \N__2689\,
            I => \N__2664\
        );

    \I__571\ : InMux
    port map (
            O => \N__2686\,
            I => \N__2664\
        );

    \I__570\ : InMux
    port map (
            O => \N__2685\,
            I => \N__2664\
        );

    \I__569\ : InMux
    port map (
            O => \N__2684\,
            I => \N__2657\
        );

    \I__568\ : InMux
    port map (
            O => \N__2683\,
            I => \N__2657\
        );

    \I__567\ : InMux
    port map (
            O => \N__2680\,
            I => \N__2657\
        );

    \I__566\ : InMux
    port map (
            O => \N__2677\,
            I => \N__2650\
        );

    \I__565\ : InMux
    port map (
            O => \N__2674\,
            I => \N__2650\
        );

    \I__564\ : InMux
    port map (
            O => \N__2671\,
            I => \N__2650\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__2664\,
            I => \greeter.M_count_qZ0Z_3\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__2657\,
            I => \greeter.M_count_qZ0Z_3\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__2650\,
            I => \greeter.M_count_qZ0Z_3\
        );

    \I__560\ : InMux
    port map (
            O => \N__2643\,
            I => \N__2632\
        );

    \I__559\ : InMux
    port map (
            O => \N__2642\,
            I => \N__2627\
        );

    \I__558\ : InMux
    port map (
            O => \N__2641\,
            I => \N__2627\
        );

    \I__557\ : InMux
    port map (
            O => \N__2640\,
            I => \N__2620\
        );

    \I__556\ : InMux
    port map (
            O => \N__2639\,
            I => \N__2620\
        );

    \I__555\ : InMux
    port map (
            O => \N__2638\,
            I => \N__2620\
        );

    \I__554\ : InMux
    port map (
            O => \N__2637\,
            I => \N__2613\
        );

    \I__553\ : InMux
    port map (
            O => \N__2636\,
            I => \N__2613\
        );

    \I__552\ : InMux
    port map (
            O => \N__2635\,
            I => \N__2613\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__2632\,
            I => \greeter.M_count_qZ0Z_0\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__2627\,
            I => \greeter.M_count_qZ0Z_0\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__2620\,
            I => \greeter.M_count_qZ0Z_0\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__2613\,
            I => \greeter.M_count_qZ0Z_0\
        );

    \I__547\ : InMux
    port map (
            O => \N__2604\,
            I => \N__2601\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__2601\,
            I => \greeter.un1_M_state_d_0_sqmuxa_1_0_a2_0_0\
        );

    \I__545\ : InMux
    port map (
            O => \N__2598\,
            I => \N__2595\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__2595\,
            I => \N__2592\
        );

    \I__543\ : Odrv12
    port map (
            O => \N__2592\,
            I => usb_rx_c
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__2589\,
            I => \N__2585\
        );

    \I__541\ : InMux
    port map (
            O => \N__2588\,
            I => \N__2581\
        );

    \I__540\ : InMux
    port map (
            O => \N__2585\,
            I => \N__2578\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__2584\,
            I => \N__2575\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__2581\,
            I => \N__2572\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__2578\,
            I => \N__2569\
        );

    \I__536\ : InMux
    port map (
            O => \N__2575\,
            I => \N__2566\
        );

    \I__535\ : Span4Mux_h
    port map (
            O => \N__2572\,
            I => \N__2563\
        );

    \I__534\ : Span4Mux_v
    port map (
            O => \N__2569\,
            I => \N__2558\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__2566\,
            I => \N__2558\
        );

    \I__532\ : Odrv4
    port map (
            O => \N__2563\,
            I => \uart_rx.M_rxd_qZ0\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__2558\,
            I => \uart_rx.M_rxd_qZ0\
        );

    \I__530\ : ClkMux
    port map (
            O => \N__2553\,
            I => \N__2508\
        );

    \I__529\ : ClkMux
    port map (
            O => \N__2552\,
            I => \N__2508\
        );

    \I__528\ : ClkMux
    port map (
            O => \N__2551\,
            I => \N__2508\
        );

    \I__527\ : ClkMux
    port map (
            O => \N__2550\,
            I => \N__2508\
        );

    \I__526\ : ClkMux
    port map (
            O => \N__2549\,
            I => \N__2508\
        );

    \I__525\ : ClkMux
    port map (
            O => \N__2548\,
            I => \N__2508\
        );

    \I__524\ : ClkMux
    port map (
            O => \N__2547\,
            I => \N__2508\
        );

    \I__523\ : ClkMux
    port map (
            O => \N__2546\,
            I => \N__2508\
        );

    \I__522\ : ClkMux
    port map (
            O => \N__2545\,
            I => \N__2508\
        );

    \I__521\ : ClkMux
    port map (
            O => \N__2544\,
            I => \N__2508\
        );

    \I__520\ : ClkMux
    port map (
            O => \N__2543\,
            I => \N__2508\
        );

    \I__519\ : ClkMux
    port map (
            O => \N__2542\,
            I => \N__2508\
        );

    \I__518\ : ClkMux
    port map (
            O => \N__2541\,
            I => \N__2508\
        );

    \I__517\ : ClkMux
    port map (
            O => \N__2540\,
            I => \N__2508\
        );

    \I__516\ : ClkMux
    port map (
            O => \N__2539\,
            I => \N__2508\
        );

    \I__515\ : GlobalMux
    port map (
            O => \N__2508\,
            I => \N__2505\
        );

    \I__514\ : gio2CtrlBuf
    port map (
            O => \N__2505\,
            I => clk_c_g
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__2502\,
            I => \M_greeter_tx_data_4_cascade_\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__2499\,
            I => \N__2495\
        );

    \I__511\ : InMux
    port map (
            O => \N__2498\,
            I => \N__2492\
        );

    \I__510\ : InMux
    port map (
            O => \N__2495\,
            I => \N__2489\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__2492\,
            I => \uart_tx.M_savedData_qZ0Z_4\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__2489\,
            I => \uart_tx.M_savedData_qZ0Z_4\
        );

    \I__507\ : CascadeMux
    port map (
            O => \N__2484\,
            I => \N__2480\
        );

    \I__506\ : InMux
    port map (
            O => \N__2483\,
            I => \N__2477\
        );

    \I__505\ : InMux
    port map (
            O => \N__2480\,
            I => \N__2474\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__2477\,
            I => \M_uart_rx_data_7\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__2474\,
            I => \M_uart_rx_data_7\
        );

    \I__502\ : InMux
    port map (
            O => \N__2469\,
            I => \N__2465\
        );

    \I__501\ : InMux
    port map (
            O => \N__2468\,
            I => \N__2462\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__2465\,
            I => \M_uart_rx_data_6\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__2462\,
            I => \M_uart_rx_data_6\
        );

    \I__498\ : InMux
    port map (
            O => \N__2457\,
            I => \N__2454\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__2454\,
            I => \M_uart_rx_data_0\
        );

    \I__496\ : InMux
    port map (
            O => \N__2451\,
            I => \N__2447\
        );

    \I__495\ : InMux
    port map (
            O => \N__2450\,
            I => \N__2444\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__2447\,
            I => \M_uart_rx_data_2\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__2444\,
            I => \M_uart_rx_data_2\
        );

    \I__492\ : InMux
    port map (
            O => \N__2439\,
            I => \N__2435\
        );

    \I__491\ : InMux
    port map (
            O => \N__2438\,
            I => \N__2432\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__2435\,
            I => \M_uart_rx_data_1\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__2432\,
            I => \M_uart_rx_data_1\
        );

    \I__488\ : InMux
    port map (
            O => \N__2427\,
            I => \N__2423\
        );

    \I__487\ : InMux
    port map (
            O => \N__2426\,
            I => \N__2420\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__2423\,
            I => \M_uart_rx_data_5\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__2420\,
            I => \M_uart_rx_data_5\
        );

    \I__484\ : CascadeMux
    port map (
            O => \N__2415\,
            I => \N_35_cascade_\
        );

    \I__483\ : InMux
    port map (
            O => \N__2412\,
            I => \N__2408\
        );

    \I__482\ : InMux
    port map (
            O => \N__2411\,
            I => \N__2405\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2408\,
            I => \uart_tx.M_savedData_qZ0Z_6\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__2405\,
            I => \uart_tx.M_savedData_qZ0Z_6\
        );

    \I__479\ : CascadeMux
    port map (
            O => \N__2400\,
            I => \N_41_cascade_\
        );

    \I__478\ : InMux
    port map (
            O => \N__2397\,
            I => \N__2393\
        );

    \I__477\ : InMux
    port map (
            O => \N__2396\,
            I => \N__2390\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__2393\,
            I => \N__2385\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__2390\,
            I => \N__2385\
        );

    \I__474\ : Odrv4
    port map (
            O => \N__2385\,
            I => \uart_tx.M_savedData_qZ0Z_2\
        );

    \I__473\ : InMux
    port map (
            O => \N__2382\,
            I => \greeter.un1_M_count_q_1_cry_0\
        );

    \I__472\ : InMux
    port map (
            O => \N__2379\,
            I => \greeter.un1_M_count_q_1_cry_1\
        );

    \I__471\ : InMux
    port map (
            O => \N__2376\,
            I => \greeter.un1_M_count_q_1_cry_2\
        );

    \I__470\ : InMux
    port map (
            O => \N__2373\,
            I => \N__2370\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__2370\,
            I => m14_0
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__2367\,
            I => \uart_rx.M_state_q_37_d_cascade_\
        );

    \I__467\ : InMux
    port map (
            O => \N__2364\,
            I => \N__2355\
        );

    \I__466\ : InMux
    port map (
            O => \N__2363\,
            I => \N__2355\
        );

    \I__465\ : InMux
    port map (
            O => \N__2362\,
            I => \N__2355\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2355\,
            I => \uart_rx.M_bitCtr_q_RNI578A4Z0Z_0\
        );

    \I__463\ : CascadeMux
    port map (
            O => \N__2352\,
            I => \N__2348\
        );

    \I__462\ : InMux
    port map (
            O => \N__2351\,
            I => \N__2339\
        );

    \I__461\ : InMux
    port map (
            O => \N__2348\,
            I => \N__2339\
        );

    \I__460\ : InMux
    port map (
            O => \N__2347\,
            I => \N__2339\
        );

    \I__459\ : InMux
    port map (
            O => \N__2346\,
            I => \N__2336\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__2339\,
            I => \uart_rx.M_bitCtr_qZ0Z_1\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__2336\,
            I => \uart_rx.M_bitCtr_qZ0Z_1\
        );

    \I__456\ : InMux
    port map (
            O => \N__2331\,
            I => \N__2325\
        );

    \I__455\ : InMux
    port map (
            O => \N__2330\,
            I => \N__2322\
        );

    \I__454\ : InMux
    port map (
            O => \N__2329\,
            I => \N__2319\
        );

    \I__453\ : InMux
    port map (
            O => \N__2328\,
            I => \N__2316\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__2325\,
            I => \uart_rx.M_ctr_q_RNILBSE3Z0Z_6\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__2322\,
            I => \uart_rx.M_ctr_q_RNILBSE3Z0Z_6\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2319\,
            I => \uart_rx.M_ctr_q_RNILBSE3Z0Z_6\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2316\,
            I => \uart_rx.M_ctr_q_RNILBSE3Z0Z_6\
        );

    \I__448\ : InMux
    port map (
            O => \N__2307\,
            I => \N__2303\
        );

    \I__447\ : InMux
    port map (
            O => \N__2306\,
            I => \N__2300\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__2303\,
            I => \uart_rx.M_bitCtr_qZ0Z_0\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__2300\,
            I => \uart_rx.M_bitCtr_qZ0Z_0\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__2295\,
            I => \greeter.M_state_q_0_cascade_\
        );

    \I__443\ : InMux
    port map (
            O => \N__2292\,
            I => \N__2289\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__2289\,
            I => \N__2286\
        );

    \I__441\ : Odrv4
    port map (
            O => \N__2286\,
            I => \greeter.M_state_d_0_sqmuxa_1_7\
        );

    \I__440\ : CascadeMux
    port map (
            O => \N__2283\,
            I => \N__2280\
        );

    \I__439\ : InMux
    port map (
            O => \N__2280\,
            I => \N__2277\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2277\,
            I => \M_uart_rx_new_data_0\
        );

    \I__437\ : InMux
    port map (
            O => \N__2274\,
            I => \N__2271\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2271\,
            I => \greeter.M_state_d_0_sqmuxa_1_6\
        );

    \I__435\ : InMux
    port map (
            O => \N__2268\,
            I => \N__2261\
        );

    \I__434\ : InMux
    port map (
            O => \N__2267\,
            I => \N__2258\
        );

    \I__433\ : InMux
    port map (
            O => \N__2266\,
            I => \N__2255\
        );

    \I__432\ : InMux
    port map (
            O => \N__2265\,
            I => \N__2250\
        );

    \I__431\ : InMux
    port map (
            O => \N__2264\,
            I => \N__2250\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2261\,
            I => \uart_tx.M_bitCtr_qZ0Z_2\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2258\,
            I => \uart_tx.M_bitCtr_qZ0Z_2\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2255\,
            I => \uart_tx.M_bitCtr_qZ0Z_2\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2250\,
            I => \uart_tx.M_bitCtr_qZ0Z_2\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__2241\,
            I => \N__2238\
        );

    \I__425\ : InMux
    port map (
            O => \N__2238\,
            I => \N__2235\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__2235\,
            I => \uart_tx.N_65\
        );

    \I__423\ : CascadeMux
    port map (
            O => \N__2232\,
            I => \N__2229\
        );

    \I__422\ : InMux
    port map (
            O => \N__2229\,
            I => \N__2223\
        );

    \I__421\ : CascadeMux
    port map (
            O => \N__2228\,
            I => \N__2220\
        );

    \I__420\ : InMux
    port map (
            O => \N__2227\,
            I => \N__2217\
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__2226\,
            I => \N__2213\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__2223\,
            I => \N__2209\
        );

    \I__417\ : InMux
    port map (
            O => \N__2220\,
            I => \N__2204\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2217\,
            I => \N__2201\
        );

    \I__415\ : InMux
    port map (
            O => \N__2216\,
            I => \N__2198\
        );

    \I__414\ : InMux
    port map (
            O => \N__2213\,
            I => \N__2193\
        );

    \I__413\ : InMux
    port map (
            O => \N__2212\,
            I => \N__2193\
        );

    \I__412\ : Span4Mux_v
    port map (
            O => \N__2209\,
            I => \N__2190\
        );

    \I__411\ : InMux
    port map (
            O => \N__2208\,
            I => \N__2185\
        );

    \I__410\ : InMux
    port map (
            O => \N__2207\,
            I => \N__2185\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2204\,
            I => \uart_rx.M_state_qZ0Z_1\
        );

    \I__408\ : Odrv12
    port map (
            O => \N__2201\,
            I => \uart_rx.M_state_qZ0Z_1\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2198\,
            I => \uart_rx.M_state_qZ0Z_1\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2193\,
            I => \uart_rx.M_state_qZ0Z_1\
        );

    \I__405\ : Odrv4
    port map (
            O => \N__2190\,
            I => \uart_rx.M_state_qZ0Z_1\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__2185\,
            I => \uart_rx.M_state_qZ0Z_1\
        );

    \I__403\ : InMux
    port map (
            O => \N__2172\,
            I => \N__2166\
        );

    \I__402\ : InMux
    port map (
            O => \N__2171\,
            I => \N__2163\
        );

    \I__401\ : InMux
    port map (
            O => \N__2170\,
            I => \N__2160\
        );

    \I__400\ : InMux
    port map (
            O => \N__2169\,
            I => \N__2157\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2166\,
            I => \uart_rx.m19_0_o2\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2163\,
            I => \uart_rx.m19_0_o2\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2160\,
            I => \uart_rx.m19_0_o2\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2157\,
            I => \uart_rx.m19_0_o2\
        );

    \I__395\ : InMux
    port map (
            O => \N__2148\,
            I => \N__2144\
        );

    \I__394\ : InMux
    port map (
            O => \N__2147\,
            I => \N__2141\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2144\,
            I => \N__2135\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2141\,
            I => \N__2132\
        );

    \I__391\ : InMux
    port map (
            O => \N__2140\,
            I => \N__2129\
        );

    \I__390\ : InMux
    port map (
            O => \N__2139\,
            I => \N__2124\
        );

    \I__389\ : InMux
    port map (
            O => \N__2138\,
            I => \N__2124\
        );

    \I__388\ : Span4Mux_s1_v
    port map (
            O => \N__2135\,
            I => \N__2117\
        );

    \I__387\ : Span4Mux_v
    port map (
            O => \N__2132\,
            I => \N__2117\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2129\,
            I => \N__2117\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2124\,
            I => \N__2114\
        );

    \I__384\ : Odrv4
    port map (
            O => \N__2117\,
            I => \M_reset_cond_out_0\
        );

    \I__383\ : Odrv4
    port map (
            O => \N__2114\,
            I => \M_reset_cond_out_0\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__2109\,
            I => \uart_rx.m19_0_0_cascade_\
        );

    \I__381\ : InMux
    port map (
            O => \N__2106\,
            I => \N__2103\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2103\,
            I => \uart_rx.M_state_d_0_sqmuxa_1\
        );

    \I__379\ : InMux
    port map (
            O => \N__2100\,
            I => \N__2096\
        );

    \I__378\ : InMux
    port map (
            O => \N__2099\,
            I => \N__2087\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2096\,
            I => \N__2084\
        );

    \I__376\ : InMux
    port map (
            O => \N__2095\,
            I => \N__2081\
        );

    \I__375\ : InMux
    port map (
            O => \N__2094\,
            I => \N__2076\
        );

    \I__374\ : InMux
    port map (
            O => \N__2093\,
            I => \N__2076\
        );

    \I__373\ : InMux
    port map (
            O => \N__2092\,
            I => \N__2073\
        );

    \I__372\ : InMux
    port map (
            O => \N__2091\,
            I => \N__2070\
        );

    \I__371\ : InMux
    port map (
            O => \N__2090\,
            I => \N__2067\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2087\,
            I => \N__2062\
        );

    \I__369\ : Span4Mux_s2_v
    port map (
            O => \N__2084\,
            I => \N__2062\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2081\,
            I => \N__2057\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2076\,
            I => \N__2057\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2073\,
            I => \uart_rx.M_state_qZ0Z_0\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2070\,
            I => \uart_rx.M_state_qZ0Z_0\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2067\,
            I => \uart_rx.M_state_qZ0Z_0\
        );

    \I__363\ : Odrv4
    port map (
            O => \N__2062\,
            I => \uart_rx.M_state_qZ0Z_0\
        );

    \I__362\ : Odrv4
    port map (
            O => \N__2057\,
            I => \uart_rx.M_state_qZ0Z_0\
        );

    \I__361\ : InMux
    port map (
            O => \N__2046\,
            I => \N__2043\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2043\,
            I => \M_greeter_tx_data_0\
        );

    \I__359\ : InMux
    port map (
            O => \N__2040\,
            I => \N__2029\
        );

    \I__358\ : InMux
    port map (
            O => \N__2039\,
            I => \N__2029\
        );

    \I__357\ : InMux
    port map (
            O => \N__2038\,
            I => \N__2026\
        );

    \I__356\ : InMux
    port map (
            O => \N__2037\,
            I => \N__2021\
        );

    \I__355\ : InMux
    port map (
            O => \N__2036\,
            I => \N__2021\
        );

    \I__354\ : InMux
    port map (
            O => \N__2035\,
            I => \N__2016\
        );

    \I__353\ : InMux
    port map (
            O => \N__2034\,
            I => \N__2016\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2029\,
            I => \uart_tx.N_183_0\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2026\,
            I => \uart_tx.N_183_0\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2021\,
            I => \uart_tx.N_183_0\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2016\,
            I => \uart_tx.N_183_0\
        );

    \I__348\ : CascadeMux
    port map (
            O => \N__2007\,
            I => \N__2004\
        );

    \I__347\ : InMux
    port map (
            O => \N__2004\,
            I => \N__1999\
        );

    \I__346\ : CascadeMux
    port map (
            O => \N__2003\,
            I => \N__1995\
        );

    \I__345\ : CascadeMux
    port map (
            O => \N__2002\,
            I => \N__1992\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__1999\,
            I => \N__1989\
        );

    \I__343\ : InMux
    port map (
            O => \N__1998\,
            I => \N__1986\
        );

    \I__342\ : InMux
    port map (
            O => \N__1995\,
            I => \N__1981\
        );

    \I__341\ : InMux
    port map (
            O => \N__1992\,
            I => \N__1981\
        );

    \I__340\ : Span4Mux_h
    port map (
            O => \N__1989\,
            I => \N__1976\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__1986\,
            I => \N__1976\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__1981\,
            I => \uart_tx.N_52_i\
        );

    \I__337\ : Odrv4
    port map (
            O => \N__1976\,
            I => \uart_tx.N_52_i\
        );

    \I__336\ : InMux
    port map (
            O => \N__1971\,
            I => \N__1968\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__1968\,
            I => \uart_tx.M_ctr_q_RNO_0Z0Z_5\
        );

    \I__334\ : InMux
    port map (
            O => \N__1965\,
            I => \N__1961\
        );

    \I__333\ : InMux
    port map (
            O => \N__1964\,
            I => \N__1958\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__1961\,
            I => \N__1955\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__1958\,
            I => \uart_tx.M_ctr_qZ0Z_5\
        );

    \I__330\ : Odrv4
    port map (
            O => \N__1955\,
            I => \uart_tx.M_ctr_qZ0Z_5\
        );

    \I__329\ : CascadeMux
    port map (
            O => \N__1950\,
            I => \greeter.M_state_d_0_sqmuxa_1_5_cascade_\
        );

    \I__328\ : CascadeMux
    port map (
            O => \N__1947\,
            I => \uart_rx.M_state_q_ns_1_cascade_\
        );

    \I__327\ : InMux
    port map (
            O => \N__1944\,
            I => \N__1937\
        );

    \I__326\ : InMux
    port map (
            O => \N__1943\,
            I => \N__1937\
        );

    \I__325\ : InMux
    port map (
            O => \N__1942\,
            I => \N__1934\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__1937\,
            I => \uart_rx.M_bitCtr_qZ0Z_2\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__1934\,
            I => \uart_rx.M_bitCtr_qZ0Z_2\
        );

    \I__322\ : InMux
    port map (
            O => \N__1929\,
            I => \N__1926\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__1926\,
            I => \uart_rx.M_state_q_37_d\
        );

    \I__320\ : InMux
    port map (
            O => \N__1923\,
            I => \N__1917\
        );

    \I__319\ : InMux
    port map (
            O => \N__1922\,
            I => \N__1917\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__1917\,
            I => \uart_tx.M_savedData_qZ0Z_0\
        );

    \I__317\ : CascadeMux
    port map (
            O => \N__1914\,
            I => \uart_tx.M_txReg_d_3_3_i_m4_ns_1_cascade_\
        );

    \I__316\ : InMux
    port map (
            O => \N__1911\,
            I => \N__1908\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__1908\,
            I => \uart_tx.N_66\
        );

    \I__314\ : CascadeMux
    port map (
            O => \N__1905\,
            I => \N__1900\
        );

    \I__313\ : CascadeMux
    port map (
            O => \N__1904\,
            I => \N__1897\
        );

    \I__312\ : CascadeMux
    port map (
            O => \N__1903\,
            I => \N__1891\
        );

    \I__311\ : InMux
    port map (
            O => \N__1900\,
            I => \N__1887\
        );

    \I__310\ : InMux
    port map (
            O => \N__1897\,
            I => \N__1882\
        );

    \I__309\ : InMux
    port map (
            O => \N__1896\,
            I => \N__1882\
        );

    \I__308\ : InMux
    port map (
            O => \N__1895\,
            I => \N__1873\
        );

    \I__307\ : InMux
    port map (
            O => \N__1894\,
            I => \N__1873\
        );

    \I__306\ : InMux
    port map (
            O => \N__1891\,
            I => \N__1873\
        );

    \I__305\ : InMux
    port map (
            O => \N__1890\,
            I => \N__1873\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__1887\,
            I => \uart_tx.M_state_qZ0Z_0\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__1882\,
            I => \uart_tx.M_state_qZ0Z_0\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__1873\,
            I => \uart_tx.M_state_qZ0Z_0\
        );

    \I__301\ : InMux
    port map (
            O => \N__1866\,
            I => \N__1863\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__1863\,
            I => \uart_tx.SUM_i_i_o4_1_1\
        );

    \I__299\ : CascadeMux
    port map (
            O => \N__1860\,
            I => \uart_tx.SUM_i_i_o4_1_1_cascade_\
        );

    \I__298\ : InMux
    port map (
            O => \N__1857\,
            I => \N__1854\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__1854\,
            I => \N__1848\
        );

    \I__296\ : InMux
    port map (
            O => \N__1853\,
            I => \N__1845\
        );

    \I__295\ : InMux
    port map (
            O => \N__1852\,
            I => \N__1840\
        );

    \I__294\ : InMux
    port map (
            O => \N__1851\,
            I => \N__1840\
        );

    \I__293\ : Odrv4
    port map (
            O => \N__1848\,
            I => \uart_tx.M_bitCtr_qZ0Z_0\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__1845\,
            I => \uart_tx.M_bitCtr_qZ0Z_0\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__1840\,
            I => \uart_tx.M_bitCtr_qZ0Z_0\
        );

    \I__290\ : CascadeMux
    port map (
            O => \N__1833\,
            I => \N__1829\
        );

    \I__289\ : InMux
    port map (
            O => \N__1832\,
            I => \N__1826\
        );

    \I__288\ : InMux
    port map (
            O => \N__1829\,
            I => \N__1816\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__1826\,
            I => \N__1813\
        );

    \I__286\ : InMux
    port map (
            O => \N__1825\,
            I => \N__1810\
        );

    \I__285\ : InMux
    port map (
            O => \N__1824\,
            I => \N__1805\
        );

    \I__284\ : InMux
    port map (
            O => \N__1823\,
            I => \N__1805\
        );

    \I__283\ : InMux
    port map (
            O => \N__1822\,
            I => \N__1802\
        );

    \I__282\ : InMux
    port map (
            O => \N__1821\,
            I => \N__1795\
        );

    \I__281\ : InMux
    port map (
            O => \N__1820\,
            I => \N__1795\
        );

    \I__280\ : InMux
    port map (
            O => \N__1819\,
            I => \N__1795\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__1816\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__278\ : Odrv4
    port map (
            O => \N__1813\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__1810\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__1805\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__1802\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__1795\,
            I => \uart_tx.M_state_qZ0Z_1\
        );

    \I__273\ : InMux
    port map (
            O => \N__1782\,
            I => \N__1776\
        );

    \I__272\ : InMux
    port map (
            O => \N__1781\,
            I => \N__1776\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__1776\,
            I => \uart_tx.M_savedData_qZ0Z_3\
        );

    \I__270\ : CascadeMux
    port map (
            O => \N__1773\,
            I => \uart_tx.M_txReg_d_0_iv_0_a2_1_1_cascade_\
        );

    \I__269\ : InMux
    port map (
            O => \N__1770\,
            I => \N__1767\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__1767\,
            I => \N__1759\
        );

    \I__267\ : InMux
    port map (
            O => \N__1766\,
            I => \N__1756\
        );

    \I__266\ : InMux
    port map (
            O => \N__1765\,
            I => \N__1753\
        );

    \I__265\ : InMux
    port map (
            O => \N__1764\,
            I => \N__1746\
        );

    \I__264\ : InMux
    port map (
            O => \N__1763\,
            I => \N__1746\
        );

    \I__263\ : InMux
    port map (
            O => \N__1762\,
            I => \N__1746\
        );

    \I__262\ : Odrv4
    port map (
            O => \N__1759\,
            I => \uart_tx.M_bitCtr_qZ0Z_1\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__1756\,
            I => \uart_tx.M_bitCtr_qZ0Z_1\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__1753\,
            I => \uart_tx.M_bitCtr_qZ0Z_1\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__1746\,
            I => \uart_tx.M_bitCtr_qZ0Z_1\
        );

    \I__258\ : InMux
    port map (
            O => \N__1737\,
            I => \N__1734\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__1734\,
            I => \N__1731\
        );

    \I__256\ : Odrv4
    port map (
            O => \N__1731\,
            I => \uart_tx.N_81\
        );

    \I__255\ : InMux
    port map (
            O => \N__1728\,
            I => \N__1725\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__1725\,
            I => \uart_tx.M_ctr_q_RNO_0Z0Z_2\
        );

    \I__253\ : InMux
    port map (
            O => \N__1722\,
            I => \N__1718\
        );

    \I__252\ : InMux
    port map (
            O => \N__1721\,
            I => \N__1715\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__1718\,
            I => \uart_tx.M_ctr_qZ0Z_2\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__1715\,
            I => \uart_tx.M_ctr_qZ0Z_2\
        );

    \I__249\ : CascadeMux
    port map (
            O => \N__1710\,
            I => \uart_rx.M_bitCtr_q_RNI578A4Z0Z_0_cascade_\
        );

    \I__248\ : InMux
    port map (
            O => \N__1707\,
            I => \N__1702\
        );

    \I__247\ : InMux
    port map (
            O => \N__1706\,
            I => \N__1699\
        );

    \I__246\ : InMux
    port map (
            O => \N__1705\,
            I => \N__1696\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__1702\,
            I => \uart_rx.M_ctr_qZ0Z_3\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__1699\,
            I => \uart_rx.M_ctr_qZ0Z_3\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__1696\,
            I => \uart_rx.M_ctr_qZ0Z_3\
        );

    \I__242\ : InMux
    port map (
            O => \N__1689\,
            I => \N__1682\
        );

    \I__241\ : InMux
    port map (
            O => \N__1688\,
            I => \N__1682\
        );

    \I__240\ : InMux
    port map (
            O => \N__1687\,
            I => \N__1679\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__1682\,
            I => \uart_rx.M_ctr_qZ0Z_5\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__1679\,
            I => \uart_rx.M_ctr_qZ0Z_5\
        );

    \I__237\ : CascadeMux
    port map (
            O => \N__1674\,
            I => \N__1671\
        );

    \I__236\ : InMux
    port map (
            O => \N__1671\,
            I => \N__1665\
        );

    \I__235\ : InMux
    port map (
            O => \N__1670\,
            I => \N__1660\
        );

    \I__234\ : InMux
    port map (
            O => \N__1669\,
            I => \N__1660\
        );

    \I__233\ : InMux
    port map (
            O => \N__1668\,
            I => \N__1657\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__1665\,
            I => \N__1654\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__1660\,
            I => \uart_rx.M_ctr_qZ0Z_2\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__1657\,
            I => \uart_rx.M_ctr_qZ0Z_2\
        );

    \I__229\ : Odrv4
    port map (
            O => \N__1654\,
            I => \uart_rx.M_ctr_qZ0Z_2\
        );

    \I__228\ : InMux
    port map (
            O => \N__1647\,
            I => \N__1642\
        );

    \I__227\ : InMux
    port map (
            O => \N__1646\,
            I => \N__1637\
        );

    \I__226\ : InMux
    port map (
            O => \N__1645\,
            I => \N__1637\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__1642\,
            I => \uart_rx.M_ctr_qZ0Z_1\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__1637\,
            I => \uart_rx.M_ctr_qZ0Z_1\
        );

    \I__223\ : InMux
    port map (
            O => \N__1632\,
            I => \N__1629\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__1629\,
            I => \uart_rx.M_ctr_q_RNIBJBV1Z0Z_1\
        );

    \I__221\ : CascadeMux
    port map (
            O => \N__1626\,
            I => \N__1623\
        );

    \I__220\ : InMux
    port map (
            O => \N__1623\,
            I => \N__1619\
        );

    \I__219\ : CascadeMux
    port map (
            O => \N__1622\,
            I => \N__1616\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1619\,
            I => \N__1612\
        );

    \I__217\ : InMux
    port map (
            O => \N__1616\,
            I => \N__1607\
        );

    \I__216\ : InMux
    port map (
            O => \N__1615\,
            I => \N__1607\
        );

    \I__215\ : Odrv4
    port map (
            O => \N__1612\,
            I => \uart_rx.M_ctr_qZ0Z_6\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__1607\,
            I => \uart_rx.M_ctr_qZ0Z_6\
        );

    \I__213\ : CascadeMux
    port map (
            O => \N__1602\,
            I => \N__1599\
        );

    \I__212\ : InMux
    port map (
            O => \N__1599\,
            I => \N__1593\
        );

    \I__211\ : InMux
    port map (
            O => \N__1598\,
            I => \N__1590\
        );

    \I__210\ : InMux
    port map (
            O => \N__1597\,
            I => \N__1587\
        );

    \I__209\ : InMux
    port map (
            O => \N__1596\,
            I => \N__1584\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__1593\,
            I => \uart_rx.M_ctr_qZ0Z_4\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__1590\,
            I => \uart_rx.M_ctr_qZ0Z_4\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__1587\,
            I => \uart_rx.M_ctr_qZ0Z_4\
        );

    \I__205\ : LocalMux
    port map (
            O => \N__1584\,
            I => \uart_rx.M_ctr_qZ0Z_4\
        );

    \I__204\ : CascadeMux
    port map (
            O => \N__1575\,
            I => \uart_rx.M_ctr_q_RNIBJBV1Z0Z_1_cascade_\
        );

    \I__203\ : InMux
    port map (
            O => \N__1572\,
            I => \N__1563\
        );

    \I__202\ : InMux
    port map (
            O => \N__1571\,
            I => \N__1563\
        );

    \I__201\ : InMux
    port map (
            O => \N__1570\,
            I => \N__1556\
        );

    \I__200\ : InMux
    port map (
            O => \N__1569\,
            I => \N__1556\
        );

    \I__199\ : InMux
    port map (
            O => \N__1568\,
            I => \N__1556\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__1563\,
            I => \uart_rx.M_ctr_qZ0Z_0\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__1556\,
            I => \uart_rx.M_ctr_qZ0Z_0\
        );

    \I__196\ : CascadeMux
    port map (
            O => \N__1551\,
            I => \uart_rx.M_ctr_q_RNILBSE3Z0Z_6_cascade_\
        );

    \I__195\ : SRMux
    port map (
            O => \N__1548\,
            I => \N__1545\
        );

    \I__194\ : LocalMux
    port map (
            O => \N__1545\,
            I => \N__1542\
        );

    \I__193\ : Span4Mux_h
    port map (
            O => \N__1542\,
            I => \N__1539\
        );

    \I__192\ : Span4Mux_s1_v
    port map (
            O => \N__1539\,
            I => \N__1536\
        );

    \I__191\ : Odrv4
    port map (
            O => \N__1536\,
            I => \uart_rx.M_state_q_RNIRDQO7_0Z0Z_0\
        );

    \I__190\ : CascadeMux
    port map (
            O => \N__1533\,
            I => \uart_tx_N_187_1_cascade_\
        );

    \I__189\ : InMux
    port map (
            O => \N__1530\,
            I => \N__1526\
        );

    \I__188\ : InMux
    port map (
            O => \N__1529\,
            I => \N__1523\
        );

    \I__187\ : LocalMux
    port map (
            O => \N__1526\,
            I => \uart_tx.N_58\
        );

    \I__186\ : LocalMux
    port map (
            O => \N__1523\,
            I => \uart_tx.N_58\
        );

    \I__185\ : InMux
    port map (
            O => \N__1518\,
            I => \N__1514\
        );

    \I__184\ : InMux
    port map (
            O => \N__1517\,
            I => \N__1511\
        );

    \I__183\ : LocalMux
    port map (
            O => \N__1514\,
            I => \uart_tx.M_ctr_qZ0Z_3\
        );

    \I__182\ : LocalMux
    port map (
            O => \N__1511\,
            I => \uart_tx.M_ctr_qZ0Z_3\
        );

    \I__181\ : InMux
    port map (
            O => \N__1506\,
            I => \uart_tx.un1_M_ctr_q_3_cry_2\
        );

    \I__180\ : InMux
    port map (
            O => \N__1503\,
            I => \N__1499\
        );

    \I__179\ : InMux
    port map (
            O => \N__1502\,
            I => \N__1496\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__1499\,
            I => \uart_tx.M_ctr_qZ0Z_4\
        );

    \I__177\ : LocalMux
    port map (
            O => \N__1496\,
            I => \uart_tx.M_ctr_qZ0Z_4\
        );

    \I__176\ : InMux
    port map (
            O => \N__1491\,
            I => \uart_tx.un1_M_ctr_q_3_cry_3\
        );

    \I__175\ : InMux
    port map (
            O => \N__1488\,
            I => \uart_tx.un1_M_ctr_q_3_cry_4\
        );

    \I__174\ : InMux
    port map (
            O => \N__1485\,
            I => \uart_tx.un1_M_ctr_q_3_cry_5\
        );

    \I__173\ : CascadeMux
    port map (
            O => \N__1482\,
            I => \uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_\
        );

    \I__172\ : CascadeMux
    port map (
            O => \N__1479\,
            I => \N__1475\
        );

    \I__171\ : InMux
    port map (
            O => \N__1478\,
            I => \N__1472\
        );

    \I__170\ : InMux
    port map (
            O => \N__1475\,
            I => \N__1469\
        );

    \I__169\ : LocalMux
    port map (
            O => \N__1472\,
            I => \uart_tx.M_ctr_qZ0Z_6\
        );

    \I__168\ : LocalMux
    port map (
            O => \N__1469\,
            I => \uart_tx.M_ctr_qZ0Z_6\
        );

    \I__167\ : IoInMux
    port map (
            O => \N__1464\,
            I => \N__1461\
        );

    \I__166\ : LocalMux
    port map (
            O => \N__1461\,
            I => usb_tx_c
        );

    \I__165\ : InMux
    port map (
            O => \N__1458\,
            I => \N__1455\
        );

    \I__164\ : LocalMux
    port map (
            O => \N__1455\,
            I => \uart_tx.M_txReg_d_0_iv_0_1\
        );

    \I__163\ : CascadeMux
    port map (
            O => \N__1452\,
            I => \N__1449\
        );

    \I__162\ : InMux
    port map (
            O => \N__1449\,
            I => \N__1439\
        );

    \I__161\ : InMux
    port map (
            O => \N__1448\,
            I => \N__1439\
        );

    \I__160\ : InMux
    port map (
            O => \N__1447\,
            I => \N__1439\
        );

    \I__159\ : InMux
    port map (
            O => \N__1446\,
            I => \N__1436\
        );

    \I__158\ : LocalMux
    port map (
            O => \N__1439\,
            I => \uart_rx.un1_M_ctr_q_5_ac0_1_out\
        );

    \I__157\ : LocalMux
    port map (
            O => \N__1436\,
            I => \uart_rx.un1_M_ctr_q_5_ac0_1_out\
        );

    \I__156\ : CascadeMux
    port map (
            O => \N__1431\,
            I => \uart_tx.M_state_q_ns_0_o2_4_0_cascade_\
        );

    \I__155\ : CascadeMux
    port map (
            O => \N__1428\,
            I => \uart_tx.N_183_0_cascade_\
        );

    \I__154\ : CascadeMux
    port map (
            O => \N__1425\,
            I => \uart_tx.M_state_q_ns_0_i_0_0_0_cascade_\
        );

    \I__153\ : CascadeMux
    port map (
            O => \N__1422\,
            I => \N__1418\
        );

    \I__152\ : InMux
    port map (
            O => \N__1421\,
            I => \N__1415\
        );

    \I__151\ : InMux
    port map (
            O => \N__1418\,
            I => \N__1412\
        );

    \I__150\ : LocalMux
    port map (
            O => \N__1415\,
            I => \uart_tx.N_187_1_i\
        );

    \I__149\ : LocalMux
    port map (
            O => \N__1412\,
            I => \uart_tx.N_187_1_i\
        );

    \I__148\ : InMux
    port map (
            O => \N__1407\,
            I => \N__1403\
        );

    \I__147\ : InMux
    port map (
            O => \N__1406\,
            I => \N__1400\
        );

    \I__146\ : LocalMux
    port map (
            O => \N__1403\,
            I => \uart_tx.M_ctr_qZ0Z_0\
        );

    \I__145\ : LocalMux
    port map (
            O => \N__1400\,
            I => \uart_tx.M_ctr_qZ0Z_0\
        );

    \I__144\ : InMux
    port map (
            O => \N__1395\,
            I => \N__1391\
        );

    \I__143\ : InMux
    port map (
            O => \N__1394\,
            I => \N__1388\
        );

    \I__142\ : LocalMux
    port map (
            O => \N__1391\,
            I => \uart_tx.M_ctr_qZ0Z_1\
        );

    \I__141\ : LocalMux
    port map (
            O => \N__1388\,
            I => \uart_tx.M_ctr_qZ0Z_1\
        );

    \I__140\ : InMux
    port map (
            O => \N__1383\,
            I => \uart_tx.un1_M_ctr_q_3_cry_0\
        );

    \I__139\ : InMux
    port map (
            O => \N__1380\,
            I => \uart_tx.un1_M_ctr_q_3_cry_1\
        );

    \I__138\ : CascadeMux
    port map (
            O => \N__1377\,
            I => \uart_rx.N_102_0_cascade_\
        );

    \I__137\ : CascadeMux
    port map (
            O => \N__1374\,
            I => \N__1370\
        );

    \I__136\ : InMux
    port map (
            O => \N__1373\,
            I => \N__1365\
        );

    \I__135\ : InMux
    port map (
            O => \N__1370\,
            I => \N__1365\
        );

    \I__134\ : LocalMux
    port map (
            O => \N__1365\,
            I => \uart_rx.un1_M_ctr_q_5_ac0_7_0\
        );

    \I__133\ : InMux
    port map (
            O => \N__1362\,
            I => \N__1344\
        );

    \I__132\ : InMux
    port map (
            O => \N__1361\,
            I => \N__1344\
        );

    \I__131\ : InMux
    port map (
            O => \N__1360\,
            I => \N__1344\
        );

    \I__130\ : InMux
    port map (
            O => \N__1359\,
            I => \N__1344\
        );

    \I__129\ : InMux
    port map (
            O => \N__1358\,
            I => \N__1344\
        );

    \I__128\ : InMux
    port map (
            O => \N__1357\,
            I => \N__1344\
        );

    \I__127\ : LocalMux
    port map (
            O => \N__1344\,
            I => \uart_rx.N_102_0\
        );

    \I__126\ : InMux
    port map (
            O => \N__1341\,
            I => \N__1338\
        );

    \I__125\ : LocalMux
    port map (
            O => \N__1338\,
            I => \uart_rx.un1_M_ctr_q_5_ac0_5_s_0_0\
        );

    \I__124\ : InMux
    port map (
            O => \N__1335\,
            I => \N__1332\
        );

    \I__123\ : LocalMux
    port map (
            O => \N__1332\,
            I => \reset_cond.M_stage_qZ0Z_1\
        );

    \I__122\ : InMux
    port map (
            O => \N__1329\,
            I => \N__1326\
        );

    \I__121\ : LocalMux
    port map (
            O => \N__1326\,
            I => \reset_cond.M_stage_qZ0Z_2\
        );

    \I__120\ : InMux
    port map (
            O => \N__1323\,
            I => \N__1311\
        );

    \I__119\ : InMux
    port map (
            O => \N__1322\,
            I => \N__1311\
        );

    \I__118\ : InMux
    port map (
            O => \N__1321\,
            I => \N__1311\
        );

    \I__117\ : InMux
    port map (
            O => \N__1320\,
            I => \N__1311\
        );

    \I__116\ : LocalMux
    port map (
            O => \N__1311\,
            I => \N__1308\
        );

    \I__115\ : IoSpan4Mux
    port map (
            O => \N__1308\,
            I => \N__1305\
        );

    \I__114\ : Odrv4
    port map (
            O => \N__1305\,
            I => rst_n_c
        );

    \I__113\ : InMux
    port map (
            O => \N__1302\,
            I => \N__1299\
        );

    \I__112\ : LocalMux
    port map (
            O => \N__1299\,
            I => \reset_cond.M_stage_qZ0Z_0\
        );

    \I__111\ : CascadeMux
    port map (
            O => \N__1296\,
            I => \uart_rx.un1_M_ctr_q_5_ac0_5_s_0_0_cascade_\
        );

    \IN_MUX_bfv_21_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_4_0_\
        );

    \IN_MUX_bfv_23_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_4_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \reset_cond.M_stage_q_1_LC_20_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__1321\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1302\,
            lcout => \reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2539\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_2_LC_20_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1322\,
            in2 => \_gnd_net_\,
            in3 => \N__1335\,
            lcout => \reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2539\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_3_LC_20_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1323\,
            in2 => \_gnd_net_\,
            in3 => \N__1329\,
            lcout => \M_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2539\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_cond.M_stage_q_0_LC_20_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1320\,
            lcout => \reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2539\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_ctr_q_RNI5PLV_3_LC_21_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1706\,
            in2 => \_gnd_net_\,
            in3 => \N__1668\,
            lcout => \uart_rx.un1_M_ctr_q_5_ac0_5_s_0_0\,
            ltout => \uart_rx.un1_M_ctr_q_5_ac0_5_s_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_ctr_q_RNIAC6F2_4_LC_21_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1446\,
            in2 => \N__1296\,
            in3 => \N__1598\,
            lcout => \uart_rx.un1_M_ctr_q_5_ac0_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_ctr_q_0_LC_21_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1571\,
            in2 => \_gnd_net_\,
            in3 => \N__1357\,
            lcout => \uart_rx.M_ctr_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2540\,
            ce => 'H',
            sr => \N__1548\
        );

    \uart_rx.M_state_q_RNIRDQO7_0_LC_21_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100000001000"
        )
    port map (
            in0 => \N__2100\,
            in1 => \N__2169\,
            in2 => \N__2232\,
            in3 => \N__2329\,
            lcout => \uart_rx.N_102_0\,
            ltout => \uart_rx.N_102_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_ctr_q_1_LC_21_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1572\,
            in2 => \N__1377\,
            in3 => \N__1647\,
            lcout => \uart_rx.M_ctr_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2540\,
            ce => 'H',
            sr => \N__1548\
        );

    \uart_rx.M_ctr_q_5_LC_21_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__1360\,
            in1 => \_gnd_net_\,
            in2 => \N__1374\,
            in3 => \N__1689\,
            lcout => \uart_rx.M_ctr_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2540\,
            ce => 'H',
            sr => \N__1548\
        );

    \uart_rx.M_ctr_q_6_LC_21_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__1688\,
            in1 => \N__1373\,
            in2 => \N__1626\,
            in3 => \N__1362\,
            lcout => \uart_rx.M_ctr_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2540\,
            ce => 'H',
            sr => \N__1548\
        );

    \uart_rx.M_ctr_q_2_LC_21_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__1358\,
            in1 => \N__1447\,
            in2 => \_gnd_net_\,
            in3 => \N__1670\,
            lcout => \uart_rx.M_ctr_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2540\,
            ce => 'H',
            sr => \N__1548\
        );

    \uart_rx.M_ctr_q_3_LC_21_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__1669\,
            in1 => \N__1361\,
            in2 => \N__1452\,
            in3 => \N__1707\,
            lcout => \uart_rx.M_ctr_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2540\,
            ce => 'H',
            sr => \N__1548\
        );

    \uart_rx.M_ctr_q_4_LC_21_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__1359\,
            in1 => \N__1448\,
            in2 => \N__1602\,
            in3 => \N__1341\,
            lcout => \uart_rx.M_ctr_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2540\,
            ce => 'H',
            sr => \N__1548\
        );

    \uart_tx.M_state_q_RNILEFM_0_LC_21_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1890\,
            in2 => \_gnd_net_\,
            in3 => \N__1819\,
            lcout => \uart_tx.N_187_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_RNILEFM_0_0_LC_21_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__1820\,
            in1 => \_gnd_net_\,
            in2 => \N__1903\,
            in3 => \_gnd_net_\,
            lcout => \uart_tx.N_52_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_1_LC_21_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__2035\,
            in1 => \N__1895\,
            in2 => \N__1833\,
            in3 => \N__2139\,
            lcout => \uart_tx.M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2542\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNIOOUF1_6_LC_21_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__1965\,
            in1 => \N__1502\,
            in2 => \N__1479\,
            in3 => \N__1394\,
            lcout => OPEN,
            ltout => \uart_tx.M_state_q_ns_0_o2_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNI3KTJ2_0_LC_21_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__1517\,
            in1 => \N__1722\,
            in2 => \N__1431\,
            in3 => \N__1407\,
            lcout => \uart_tx.N_183_0\,
            ltout => \uart_tx.N_183_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_RNIR97K3_1_LC_21_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1866\,
            in2 => \N__1428\,
            in3 => \N__1765\,
            lcout => \uart_tx.N_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_RNO_0_0_LC_21_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110100"
        )
    port map (
            in0 => \N__2034\,
            in1 => \N__1894\,
            in2 => \N__2984\,
            in3 => \N__1821\,
            lcout => OPEN,
            ltout => \uart_tx.M_state_q_ns_0_i_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_0_LC_21_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010100"
        )
    port map (
            in0 => \N__2138\,
            in1 => \N__2268\,
            in2 => \N__1425\,
            in3 => \N__1530\,
            lcout => \uart_tx.M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2542\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_0_LC_21_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2870\,
            in1 => \N__1406\,
            in2 => \N__1422\,
            in3 => \N__1421\,
            lcout => \uart_tx.M_ctr_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_21_4_0_\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_0\,
            clk => \N__2544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_1_LC_21_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2874\,
            in1 => \N__1395\,
            in2 => \_gnd_net_\,
            in3 => \N__1383\,
            lcout => \uart_tx.M_ctr_qZ0Z_1\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_0\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_1\,
            clk => \N__2544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNO_0_2_LC_21_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1721\,
            in2 => \_gnd_net_\,
            in3 => \N__1380\,
            lcout => \uart_tx.M_ctr_q_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_1\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_3_LC_21_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2873\,
            in1 => \N__1518\,
            in2 => \_gnd_net_\,
            in3 => \N__1506\,
            lcout => \uart_tx.M_ctr_qZ0Z_3\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_2\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_3\,
            clk => \N__2544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_4_LC_21_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2871\,
            in1 => \N__1503\,
            in2 => \_gnd_net_\,
            in3 => \N__1491\,
            lcout => \uart_tx.M_ctr_qZ0Z_4\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_3\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_4\,
            clk => \N__2544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNO_0_5_LC_21_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1964\,
            in2 => \_gnd_net_\,
            in3 => \N__1488\,
            lcout => \uart_tx.M_ctr_q_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \uart_tx.un1_M_ctr_q_3_cry_4\,
            carryout => \uart_tx.un1_M_ctr_q_3_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_RNO_0_6_LC_21_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1478\,
            in2 => \_gnd_net_\,
            in3 => \N__1485\,
            lcout => OPEN,
            ltout => \uart_tx.M_ctr_q_RNO_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_6_LC_21_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__1998\,
            in1 => \N__2872\,
            in2 => \N__1482\,
            in3 => \N__2038\,
            lcout => \uart_tx.M_ctr_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2544\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_LC_22_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111110101111"
        )
    port map (
            in0 => \N__1737\,
            in1 => \N__1458\,
            in2 => \N__2007\,
            in3 => \N__1832\,
            lcout => usb_tx_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2541\,
            ce => 'H',
            sr => \N__2892\
        );

    \uart_tx.M_txReg_q_RNO_1_LC_22_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__1857\,
            in1 => \N__1911\,
            in2 => \N__2241\,
            in3 => \N__1770\,
            lcout => \uart_tx.M_txReg_d_0_iv_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_ctr_q_RNI1LLV_1_LC_22_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__1569\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1646\,
            lcout => \uart_rx.un1_M_ctr_q_5_ac0_1_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_state_q_ns_1_0__m19_0_o2_LC_22_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__1597\,
            in1 => \N__1570\,
            in2 => \N__1622\,
            in3 => \N__1632\,
            lcout => \uart_rx.m19_0_o2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_bitCtr_q_RNI578A4_0_LC_22_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__2090\,
            in1 => \N__2306\,
            in2 => \N__2226\,
            in3 => \N__2328\,
            lcout => \uart_rx.M_bitCtr_q_RNI578A4Z0Z_0\,
            ltout => \uart_rx.M_bitCtr_q_RNI578A4Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_state_q_ns_1_0__m19_0_a2_1_LC_22_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__2346\,
            in1 => \_gnd_net_\,
            in2 => \N__1710\,
            in3 => \N__1942\,
            lcout => \uart_rx.M_state_d_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_ctr_q_RNIBJBV1_1_LC_22_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__1705\,
            in1 => \N__1687\,
            in2 => \N__1674\,
            in3 => \N__1645\,
            lcout => \uart_rx.M_ctr_q_RNIBJBV1Z0Z_1\,
            ltout => \uart_rx.M_ctr_q_RNIBJBV1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_ctr_q_RNILBSE3_6_LC_22_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__1615\,
            in1 => \N__1596\,
            in2 => \N__1575\,
            in3 => \N__1568\,
            lcout => \uart_rx.M_ctr_q_RNILBSE3Z0Z_6\,
            ltout => \uart_rx.M_ctr_q_RNILBSE3Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_state_q_RNIRDQO7_0_0_LC_22_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101010111"
        )
    port map (
            in0 => \N__2212\,
            in1 => \N__2095\,
            in2 => \N__1551\,
            in3 => \N__2172\,
            lcout => \uart_rx.M_state_q_RNIRDQO7_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_0_LC_22_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__2046\,
            in1 => \N__2876\,
            in2 => \N__2977\,
            in3 => \N__1923\,
            lcout => \uart_tx.M_savedData_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_state_q_RNILEFM_1_0_LC_22_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1896\,
            in2 => \_gnd_net_\,
            in3 => \N__1822\,
            lcout => \uart_tx_N_187_1\,
            ltout => \uart_tx_N_187_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_2_LC_22_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__2265\,
            in1 => \_gnd_net_\,
            in2 => \N__1533\,
            in3 => \N__1529\,
            lcout => \uart_tx.M_bitCtr_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_5_LC_22_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__1922\,
            in1 => \N__2264\,
            in2 => \N__2499\,
            in3 => \N__1762\,
            lcout => OPEN,
            ltout => \uart_tx.M_txReg_d_3_3_i_m4_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_4_LC_22_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__1763\,
            in1 => \N__2411\,
            in2 => \N__1914\,
            in3 => \N__2396\,
            lcout => \uart_tx.N_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_0_LC_22_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000001000"
        )
    port map (
            in0 => \N__1824\,
            in1 => \N__2037\,
            in2 => \N__1905\,
            in3 => \N__1852\,
            lcout => \uart_tx.M_bitCtr_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_RNIMHCR_0_LC_22_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__1851\,
            in1 => \_gnd_net_\,
            in2 => \N__1904\,
            in3 => \N__1823\,
            lcout => \uart_tx.SUM_i_i_o4_1_1\,
            ltout => \uart_tx.SUM_i_i_o4_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_bitCtr_q_1_LC_22_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000100000100"
        )
    port map (
            in0 => \N__2875\,
            in1 => \N__2036\,
            in2 => \N__1860\,
            in3 => \N__1764\,
            lcout => \uart_tx.M_bitCtr_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2545\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_3_LC_22_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101011101010"
        )
    port map (
            in0 => \N__1782\,
            in1 => \N__2879\,
            in2 => \N__2985\,
            in3 => \N__2373\,
            lcout => \uart_tx.M_savedData_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_2_LC_22_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1853\,
            in2 => \_gnd_net_\,
            in3 => \N__1825\,
            lcout => OPEN,
            ltout => \uart_tx.M_txReg_d_0_iv_0_a2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_0_LC_22_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2267\,
            in1 => \N__1781\,
            in2 => \N__1773\,
            in3 => \N__1766\,
            lcout => \uart_tx.N_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_2_LC_22_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__2877\,
            in1 => \N__2039\,
            in2 => \N__2002\,
            in3 => \N__1728\,
            lcout => \uart_tx.M_ctr_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_ctr_q_5_LC_22_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__2878\,
            in1 => \N__2040\,
            in2 => \N__2003\,
            in3 => \N__1971\,
            lcout => \uart_tx.M_ctr_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2548\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.M_state_q_RNO_3_LC_23_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__2426\,
            in1 => \N__3044\,
            in2 => \N__2484\,
            in3 => \N__3032\,
            lcout => OPEN,
            ltout => \greeter.M_state_d_0_sqmuxa_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.M_state_q_RNO_1_LC_23_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__2457\,
            in1 => \_gnd_net_\,
            in2 => \N__1950\,
            in3 => \N__2939\,
            lcout => \greeter.M_state_d_0_sqmuxa_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_state_q_ns_1_0__m22_0_LC_23_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101001101110"
        )
    port map (
            in0 => \N__2208\,
            in1 => \N__2094\,
            in2 => \N__2584\,
            in3 => \N__2170\,
            lcout => OPEN,
            ltout => \uart_rx.M_state_q_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_state_q_1_LC_23_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1947\,
            in3 => \N__2148\,
            lcout => \uart_rx.M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_state_q_RNI62U94_0_LC_23_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__2207\,
            in1 => \N__2093\,
            in2 => \_gnd_net_\,
            in3 => \N__2330\,
            lcout => \uart_rx.N_25_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_bitCtr_q_2_LC_23_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100010000"
        )
    port map (
            in0 => \N__2363\,
            in1 => \N__1929\,
            in2 => \N__2352\,
            in3 => \N__1943\,
            lcout => \uart_rx.M_bitCtr_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2546\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_newData_q_LC_23_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__1944\,
            in1 => \N__2351\,
            in2 => \_gnd_net_\,
            in3 => \N__2364\,
            lcout => \M_uart_rx_new_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2546\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_state_q_RNIHM1R_0_LC_23_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2216\,
            in2 => \_gnd_net_\,
            in3 => \N__2091\,
            lcout => \uart_rx.M_state_q_37_d\,
            ltout => \uart_rx.M_state_q_37_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_bitCtr_q_1_LC_23_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2347\,
            in2 => \N__2367\,
            in3 => \N__2362\,
            lcout => \uart_rx.M_bitCtr_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2546\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_bitCtr_q_0_LC_23_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100010011000"
        )
    port map (
            in0 => \N__2092\,
            in1 => \N__2307\,
            in2 => \N__2228\,
            in3 => \N__2331\,
            lcout => \uart_rx.M_bitCtr_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2546\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.M_state_q_RNO_2_LC_23_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__2940\,
            in1 => \N__2604\,
            in2 => \_gnd_net_\,
            in3 => \N__2859\,
            lcout => OPEN,
            ltout => \greeter.M_state_q_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.M_state_q_LC_23_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010001010000"
        )
    port map (
            in0 => \N__2140\,
            in1 => \N__2274\,
            in2 => \N__2295\,
            in3 => \N__2292\,
            lcout => \greeter_M_state_q\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2546\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.M_state_q_RNO_0_LC_23_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__2468\,
            in1 => \N__2450\,
            in2 => \N__2283\,
            in3 => \N__2438\,
            lcout => \greeter.M_state_d_0_sqmuxa_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_txReg_q_RNO_3_LC_23_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__2996\,
            in1 => \N__2789\,
            in2 => \_gnd_net_\,
            in3 => \N__2266\,
            lcout => \uart_tx.N_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_state_q_ns_1_0__m19_0_0_LC_23_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001001"
        )
    port map (
            in0 => \N__2227\,
            in1 => \N__2099\,
            in2 => \N__2589\,
            in3 => \N__2171\,
            lcout => OPEN,
            ltout => \uart_rx.m19_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_state_q_0_LC_23_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010000"
        )
    port map (
            in0 => \N__2147\,
            in1 => \_gnd_net_\,
            in2 => \N__2109\,
            in3 => \N__2106\,
            lcout => \uart_rx.M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2549\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.rom.letter_1_6_0__m5_0_LC_23_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101110000100"
        )
    port map (
            in0 => \N__2725\,
            in1 => \N__2638\,
            in2 => \N__2693\,
            in3 => \N__2764\,
            lcout => \M_greeter_tx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.rom.letter_1_6_0__m23_i_LC_23_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000100000"
        )
    port map (
            in0 => \N__2640\,
            in1 => \N__2727\,
            in2 => \N__2778\,
            in3 => \N__2684\,
            lcout => OPEN,
            ltout => \N_35_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_6_LC_23_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__2960\,
            in1 => \N__2412\,
            in2 => \N__2415\,
            in3 => \N__2888\,
            lcout => \uart_tx.M_savedData_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2549\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.rom.letter_1_6_0__m12_i_LC_23_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100100100001"
        )
    port map (
            in0 => \N__2639\,
            in1 => \N__2726\,
            in2 => \N__2777\,
            in3 => \N__2683\,
            lcout => OPEN,
            ltout => \N_41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_2_LC_23_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__2959\,
            in1 => \N__2397\,
            in2 => \N__2400\,
            in3 => \N__2887\,
            lcout => \uart_tx.M_savedData_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2549\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.M_count_q_0_LC_23_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__2972\,
            in1 => \N__2643\,
            in2 => \N__2884\,
            in3 => \N__2880\,
            lcout => \greeter.M_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_23_4_0_\,
            carryout => \greeter.un1_M_count_q_1_cry_0\,
            clk => \N__2551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.M_count_q_1_LC_23_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__2975\,
            in1 => \N__2732\,
            in2 => \_gnd_net_\,
            in3 => \N__2382\,
            lcout => \greeter.M_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \greeter.un1_M_count_q_1_cry_0\,
            carryout => \greeter.un1_M_count_q_1_cry_1\,
            clk => \N__2551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.M_count_q_2_LC_23_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__2973\,
            in1 => \N__2773\,
            in2 => \_gnd_net_\,
            in3 => \N__2379\,
            lcout => \greeter.M_count_qZ1Z_2\,
            ltout => OPEN,
            carryin => \greeter.un1_M_count_q_1_cry_1\,
            carryout => \greeter.un1_M_count_q_1_cry_2\,
            clk => \N__2551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.M_count_q_3_LC_23_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__2689\,
            in1 => \N__2974\,
            in2 => \_gnd_net_\,
            in3 => \N__2376\,
            lcout => \greeter.M_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.rom.letter_1_6_0__m14_0_LC_23_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001101011000"
        )
    port map (
            in0 => \N__2771\,
            in1 => \N__2728\,
            in2 => \N__2694\,
            in3 => \N__2641\,
            lcout => m14_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.rom.letter_1_6_0__m17_0_LC_23_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000100"
        )
    port map (
            in0 => \N__2642\,
            in1 => \N__2685\,
            in2 => \N__2733\,
            in3 => \N__2772\,
            lcout => OPEN,
            ltout => \M_greeter_tx_data_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_4_LC_23_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__2976\,
            in1 => \N__2858\,
            in2 => \N__2502\,
            in3 => \N__2498\,
            lcout => \uart_tx.M_savedData_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2551\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_savedData_q_6_LC_24_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2483\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_uart_rx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2547\,
            ce => \N__3017\,
            sr => \_gnd_net_\
        );

    \uart_rx.M_savedData_q_7_LC_24_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2588\,
            lcout => \M_uart_rx_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2550\,
            ce => \N__3021\,
            sr => \_gnd_net_\
        );

    \uart_rx.M_savedData_q_2_LC_24_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3033\,
            lcout => \M_uart_rx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2550\,
            ce => \N__3021\,
            sr => \_gnd_net_\
        );

    \uart_rx.M_savedData_q_5_LC_24_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2469\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_uart_rx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2550\,
            ce => \N__3021\,
            sr => \_gnd_net_\
        );

    \uart_rx.M_savedData_q_0_LC_24_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2439\,
            lcout => \M_uart_rx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2550\,
            ce => \N__3021\,
            sr => \_gnd_net_\
        );

    \uart_rx.M_savedData_q_1_LC_24_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2451\,
            lcout => \M_uart_rx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2550\,
            ce => \N__3021\,
            sr => \_gnd_net_\
        );

    \uart_rx.M_savedData_q_4_LC_24_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2427\,
            lcout => \M_uart_rx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2550\,
            ce => \N__3021\,
            sr => \_gnd_net_\
        );

    \uart_rx.M_savedData_q_3_LC_24_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3045\,
            lcout => \M_uart_rx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2550\,
            ce => \N__3021\,
            sr => \_gnd_net_\
        );

    \greeter.rom.letter_1_6_0__m20_i_LC_24_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101001"
        )
    port map (
            in0 => \N__2775\,
            in1 => \N__2723\,
            in2 => \N__2691\,
            in3 => \N__2636\,
            lcout => OPEN,
            ltout => \N_37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_5_LC_24_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__2965\,
            in1 => \N__2997\,
            in2 => \N__3000\,
            in3 => \N__2886\,
            lcout => \uart_tx.M_savedData_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.rom.letter_1_6_0__m9_0_LC_24_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000111010"
        )
    port map (
            in0 => \N__2776\,
            in1 => \N__2724\,
            in2 => \N__2692\,
            in3 => \N__2637\,
            lcout => OPEN,
            ltout => \M_greeter_tx_data_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_tx.M_savedData_q_1_LC_24_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__2964\,
            in1 => \N__2790\,
            in2 => \N__2895\,
            in3 => \N__2885\,
            lcout => \uart_tx.M_savedData_qZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \greeter.M_state_q_RNO_4_LC_24_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2774\,
            in1 => \N__2722\,
            in2 => \N__2690\,
            in3 => \N__2635\,
            lcout => \greeter.un1_M_state_d_0_sqmuxa_1_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_rx.M_rxd_q_LC_26_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2598\,
            lcout => \uart_rx.M_rxd_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2553\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
